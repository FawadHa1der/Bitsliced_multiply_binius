module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 ;
  assign n628 = x31 & x63 ;
  assign n627 = x30 & x62 ;
  assign n632 = n628 ^ n627 ;
  assign n621 = x29 & x61 ;
  assign n620 = x28 & x60 ;
  assign n625 = n621 ^ n620 ;
  assign n646 = n632 ^ n625 ;
  assign n596 = x27 & x59 ;
  assign n595 = x26 & x58 ;
  assign n600 = n596 ^ n595 ;
  assign n589 = x25 & x57 ;
  assign n588 = x24 & x56 ;
  assign n593 = n589 ^ n588 ;
  assign n614 = n600 ^ n593 ;
  assign n695 = n646 ^ n614 ;
  assign n509 = x23 & x55 ;
  assign n508 = x22 & x54 ;
  assign n513 = n509 ^ n508 ;
  assign n502 = x21 & x53 ;
  assign n501 = x20 & x52 ;
  assign n506 = n502 ^ n501 ;
  assign n527 = n513 ^ n506 ;
  assign n477 = x19 & x51 ;
  assign n476 = x18 & x50 ;
  assign n481 = n477 ^ n476 ;
  assign n470 = x17 & x49 ;
  assign n469 = x16 & x48 ;
  assign n474 = n470 ^ n469 ;
  assign n495 = n481 ^ n474 ;
  assign n576 = n527 ^ n495 ;
  assign n849 = n695 ^ n576 ;
  assign n224 = x15 & x47 ;
  assign n223 = x14 & x46 ;
  assign n228 = n224 ^ n223 ;
  assign n217 = x13 & x45 ;
  assign n216 = x12 & x44 ;
  assign n221 = n217 ^ n216 ;
  assign n242 = n228 ^ n221 ;
  assign n192 = x11 & x43 ;
  assign n191 = x10 & x42 ;
  assign n196 = n192 ^ n191 ;
  assign n185 = x9 & x41 ;
  assign n184 = x8 & x40 ;
  assign n189 = n185 ^ n184 ;
  assign n210 = n196 ^ n189 ;
  assign n291 = n242 ^ n210 ;
  assign n105 = x7 & x39 ;
  assign n104 = x6 & x38 ;
  assign n109 = n105 ^ n104 ;
  assign n98 = x5 & x37 ;
  assign n97 = x4 & x36 ;
  assign n102 = n98 ^ n97 ;
  assign n123 = n109 ^ n102 ;
  assign n73 = x3 & x35 ;
  assign n72 = x2 & x34 ;
  assign n77 = n73 ^ n72 ;
  assign n66 = x1 & x33 ;
  assign n65 = x0 & x32 ;
  assign n70 = n66 ^ n65 ;
  assign n91 = n77 ^ n70 ;
  assign n172 = n123 ^ n91 ;
  assign n445 = n291 ^ n172 ;
  assign n1324 = n849 ^ n445 ;
  assign n629 = x31 ^ x30 ;
  assign n630 = x63 ^ x62 ;
  assign n631 = n629 & n630 ;
  assign n633 = n631 ^ n627 ;
  assign n622 = x29 ^ x28 ;
  assign n623 = x61 ^ x60 ;
  assign n624 = n622 & n623 ;
  assign n626 = n624 ^ n620 ;
  assign n647 = n633 ^ n626 ;
  assign n597 = x27 ^ x26 ;
  assign n598 = x59 ^ x58 ;
  assign n599 = n597 & n598 ;
  assign n601 = n599 ^ n595 ;
  assign n590 = x25 ^ x24 ;
  assign n591 = x57 ^ x56 ;
  assign n592 = n590 & n591 ;
  assign n594 = n592 ^ n588 ;
  assign n615 = n601 ^ n594 ;
  assign n696 = n647 ^ n615 ;
  assign n510 = x23 ^ x22 ;
  assign n511 = x55 ^ x54 ;
  assign n512 = n510 & n511 ;
  assign n514 = n512 ^ n508 ;
  assign n503 = x21 ^ x20 ;
  assign n504 = x53 ^ x52 ;
  assign n505 = n503 & n504 ;
  assign n507 = n505 ^ n501 ;
  assign n528 = n514 ^ n507 ;
  assign n478 = x19 ^ x18 ;
  assign n479 = x51 ^ x50 ;
  assign n480 = n478 & n479 ;
  assign n482 = n480 ^ n476 ;
  assign n471 = x17 ^ x16 ;
  assign n472 = x49 ^ x48 ;
  assign n473 = n471 & n472 ;
  assign n475 = n473 ^ n469 ;
  assign n496 = n482 ^ n475 ;
  assign n577 = n528 ^ n496 ;
  assign n850 = n696 ^ n577 ;
  assign n225 = x15 ^ x14 ;
  assign n226 = x47 ^ x46 ;
  assign n227 = n225 & n226 ;
  assign n229 = n227 ^ n223 ;
  assign n218 = x13 ^ x12 ;
  assign n219 = x45 ^ x44 ;
  assign n220 = n218 & n219 ;
  assign n222 = n220 ^ n216 ;
  assign n243 = n229 ^ n222 ;
  assign n193 = x11 ^ x10 ;
  assign n194 = x43 ^ x42 ;
  assign n195 = n193 & n194 ;
  assign n197 = n195 ^ n191 ;
  assign n186 = x9 ^ x8 ;
  assign n187 = x41 ^ x40 ;
  assign n188 = n186 & n187 ;
  assign n190 = n188 ^ n184 ;
  assign n211 = n197 ^ n190 ;
  assign n292 = n243 ^ n211 ;
  assign n106 = x7 ^ x6 ;
  assign n107 = x39 ^ x38 ;
  assign n108 = n106 & n107 ;
  assign n110 = n108 ^ n104 ;
  assign n99 = x5 ^ x4 ;
  assign n100 = x37 ^ x36 ;
  assign n101 = n99 & n100 ;
  assign n103 = n101 ^ n97 ;
  assign n124 = n110 ^ n103 ;
  assign n74 = x3 ^ x2 ;
  assign n75 = x35 ^ x34 ;
  assign n76 = n74 & n75 ;
  assign n78 = n76 ^ n72 ;
  assign n67 = x1 ^ x0 ;
  assign n68 = x33 ^ x32 ;
  assign n69 = n67 & n68 ;
  assign n71 = n69 ^ n65 ;
  assign n92 = n78 ^ n71 ;
  assign n173 = n124 ^ n92 ;
  assign n446 = n292 ^ n173 ;
  assign n1325 = n850 ^ n446 ;
  assign n636 = x31 ^ x29 ;
  assign n637 = x63 ^ x61 ;
  assign n640 = n636 & n637 ;
  assign n634 = x30 ^ x28 ;
  assign n635 = x62 ^ x60 ;
  assign n639 = n634 & n635 ;
  assign n644 = n640 ^ n639 ;
  assign n648 = n646 ^ n644 ;
  assign n649 = n648 ^ n633 ;
  assign n604 = x27 ^ x25 ;
  assign n605 = x59 ^ x57 ;
  assign n608 = n604 & n605 ;
  assign n602 = x26 ^ x24 ;
  assign n603 = x58 ^ x56 ;
  assign n607 = n602 & n603 ;
  assign n612 = n608 ^ n607 ;
  assign n616 = n614 ^ n612 ;
  assign n617 = n616 ^ n601 ;
  assign n697 = n649 ^ n617 ;
  assign n517 = x23 ^ x21 ;
  assign n518 = x55 ^ x53 ;
  assign n521 = n517 & n518 ;
  assign n515 = x22 ^ x20 ;
  assign n516 = x54 ^ x52 ;
  assign n520 = n515 & n516 ;
  assign n525 = n521 ^ n520 ;
  assign n529 = n527 ^ n525 ;
  assign n530 = n529 ^ n514 ;
  assign n485 = x19 ^ x17 ;
  assign n486 = x51 ^ x49 ;
  assign n489 = n485 & n486 ;
  assign n483 = x18 ^ x16 ;
  assign n484 = x50 ^ x48 ;
  assign n488 = n483 & n484 ;
  assign n493 = n489 ^ n488 ;
  assign n497 = n495 ^ n493 ;
  assign n498 = n497 ^ n482 ;
  assign n578 = n530 ^ n498 ;
  assign n851 = n697 ^ n578 ;
  assign n232 = x15 ^ x13 ;
  assign n233 = x47 ^ x45 ;
  assign n236 = n232 & n233 ;
  assign n230 = x14 ^ x12 ;
  assign n231 = x46 ^ x44 ;
  assign n235 = n230 & n231 ;
  assign n240 = n236 ^ n235 ;
  assign n244 = n242 ^ n240 ;
  assign n245 = n244 ^ n229 ;
  assign n200 = x11 ^ x9 ;
  assign n201 = x43 ^ x41 ;
  assign n204 = n200 & n201 ;
  assign n198 = x10 ^ x8 ;
  assign n199 = x42 ^ x40 ;
  assign n203 = n198 & n199 ;
  assign n208 = n204 ^ n203 ;
  assign n212 = n210 ^ n208 ;
  assign n213 = n212 ^ n197 ;
  assign n293 = n245 ^ n213 ;
  assign n113 = x7 ^ x5 ;
  assign n114 = x39 ^ x37 ;
  assign n117 = n113 & n114 ;
  assign n111 = x6 ^ x4 ;
  assign n112 = x38 ^ x36 ;
  assign n116 = n111 & n112 ;
  assign n121 = n117 ^ n116 ;
  assign n125 = n123 ^ n121 ;
  assign n126 = n125 ^ n110 ;
  assign n81 = x3 ^ x1 ;
  assign n82 = x35 ^ x33 ;
  assign n85 = n81 & n82 ;
  assign n79 = x2 ^ x0 ;
  assign n80 = x34 ^ x32 ;
  assign n84 = n79 & n80 ;
  assign n89 = n85 ^ n84 ;
  assign n93 = n91 ^ n89 ;
  assign n94 = n93 ^ n78 ;
  assign n174 = n126 ^ n94 ;
  assign n447 = n293 ^ n174 ;
  assign n1326 = n851 ^ n447 ;
  assign n641 = n636 ^ n634 ;
  assign n642 = n637 ^ n635 ;
  assign n643 = n641 & n642 ;
  assign n645 = n643 ^ n639 ;
  assign n650 = n647 ^ n645 ;
  assign n638 = n633 ^ n632 ;
  assign n651 = n650 ^ n638 ;
  assign n609 = n604 ^ n602 ;
  assign n610 = n605 ^ n603 ;
  assign n611 = n609 & n610 ;
  assign n613 = n611 ^ n607 ;
  assign n618 = n615 ^ n613 ;
  assign n606 = n601 ^ n600 ;
  assign n619 = n618 ^ n606 ;
  assign n698 = n651 ^ n619 ;
  assign n522 = n517 ^ n515 ;
  assign n523 = n518 ^ n516 ;
  assign n524 = n522 & n523 ;
  assign n526 = n524 ^ n520 ;
  assign n531 = n528 ^ n526 ;
  assign n519 = n514 ^ n513 ;
  assign n532 = n531 ^ n519 ;
  assign n490 = n485 ^ n483 ;
  assign n491 = n486 ^ n484 ;
  assign n492 = n490 & n491 ;
  assign n494 = n492 ^ n488 ;
  assign n499 = n496 ^ n494 ;
  assign n487 = n482 ^ n481 ;
  assign n500 = n499 ^ n487 ;
  assign n579 = n532 ^ n500 ;
  assign n852 = n698 ^ n579 ;
  assign n237 = n232 ^ n230 ;
  assign n238 = n233 ^ n231 ;
  assign n239 = n237 & n238 ;
  assign n241 = n239 ^ n235 ;
  assign n246 = n243 ^ n241 ;
  assign n234 = n229 ^ n228 ;
  assign n247 = n246 ^ n234 ;
  assign n205 = n200 ^ n198 ;
  assign n206 = n201 ^ n199 ;
  assign n207 = n205 & n206 ;
  assign n209 = n207 ^ n203 ;
  assign n214 = n211 ^ n209 ;
  assign n202 = n197 ^ n196 ;
  assign n215 = n214 ^ n202 ;
  assign n294 = n247 ^ n215 ;
  assign n118 = n113 ^ n111 ;
  assign n119 = n114 ^ n112 ;
  assign n120 = n118 & n119 ;
  assign n122 = n120 ^ n116 ;
  assign n127 = n124 ^ n122 ;
  assign n115 = n110 ^ n109 ;
  assign n128 = n127 ^ n115 ;
  assign n86 = n81 ^ n79 ;
  assign n87 = n82 ^ n80 ;
  assign n88 = n86 & n87 ;
  assign n90 = n88 ^ n84 ;
  assign n95 = n92 ^ n90 ;
  assign n83 = n78 ^ n77 ;
  assign n96 = n95 ^ n83 ;
  assign n175 = n128 ^ n96 ;
  assign n448 = n294 ^ n175 ;
  assign n1327 = n852 ^ n448 ;
  assign n658 = x31 ^ x27 ;
  assign n659 = x63 ^ x59 ;
  assign n671 = n658 & n659 ;
  assign n656 = x30 ^ x26 ;
  assign n657 = x62 ^ x58 ;
  assign n670 = n656 & n657 ;
  assign n675 = n671 ^ n670 ;
  assign n654 = x29 ^ x25 ;
  assign n655 = x61 ^ x57 ;
  assign n664 = n654 & n655 ;
  assign n652 = x28 ^ x24 ;
  assign n653 = x60 ^ x56 ;
  assign n663 = n652 & n653 ;
  assign n668 = n664 ^ n663 ;
  assign n689 = n675 ^ n668 ;
  assign n699 = n695 ^ n689 ;
  assign n700 = n699 ^ n649 ;
  assign n539 = x23 ^ x19 ;
  assign n540 = x55 ^ x51 ;
  assign n552 = n539 & n540 ;
  assign n537 = x22 ^ x18 ;
  assign n538 = x54 ^ x50 ;
  assign n551 = n537 & n538 ;
  assign n556 = n552 ^ n551 ;
  assign n535 = x21 ^ x17 ;
  assign n536 = x53 ^ x49 ;
  assign n545 = n535 & n536 ;
  assign n533 = x20 ^ x16 ;
  assign n534 = x52 ^ x48 ;
  assign n544 = n533 & n534 ;
  assign n549 = n545 ^ n544 ;
  assign n570 = n556 ^ n549 ;
  assign n580 = n576 ^ n570 ;
  assign n581 = n580 ^ n530 ;
  assign n853 = n700 ^ n581 ;
  assign n254 = x15 ^ x11 ;
  assign n255 = x47 ^ x43 ;
  assign n267 = n254 & n255 ;
  assign n252 = x14 ^ x10 ;
  assign n253 = x46 ^ x42 ;
  assign n266 = n252 & n253 ;
  assign n271 = n267 ^ n266 ;
  assign n250 = x13 ^ x9 ;
  assign n251 = x45 ^ x41 ;
  assign n260 = n250 & n251 ;
  assign n248 = x12 ^ x8 ;
  assign n249 = x44 ^ x40 ;
  assign n259 = n248 & n249 ;
  assign n264 = n260 ^ n259 ;
  assign n285 = n271 ^ n264 ;
  assign n295 = n291 ^ n285 ;
  assign n296 = n295 ^ n245 ;
  assign n135 = x7 ^ x3 ;
  assign n136 = x39 ^ x35 ;
  assign n148 = n135 & n136 ;
  assign n133 = x6 ^ x2 ;
  assign n134 = x38 ^ x34 ;
  assign n147 = n133 & n134 ;
  assign n152 = n148 ^ n147 ;
  assign n131 = x5 ^ x1 ;
  assign n132 = x37 ^ x33 ;
  assign n141 = n131 & n132 ;
  assign n129 = x4 ^ x0 ;
  assign n130 = x36 ^ x32 ;
  assign n140 = n129 & n130 ;
  assign n145 = n141 ^ n140 ;
  assign n166 = n152 ^ n145 ;
  assign n176 = n172 ^ n166 ;
  assign n177 = n176 ^ n126 ;
  assign n449 = n296 ^ n177 ;
  assign n1328 = n853 ^ n449 ;
  assign n672 = n658 ^ n656 ;
  assign n673 = n659 ^ n657 ;
  assign n674 = n672 & n673 ;
  assign n676 = n674 ^ n670 ;
  assign n665 = n654 ^ n652 ;
  assign n666 = n655 ^ n653 ;
  assign n667 = n665 & n666 ;
  assign n669 = n667 ^ n663 ;
  assign n690 = n676 ^ n669 ;
  assign n701 = n696 ^ n690 ;
  assign n702 = n701 ^ n651 ;
  assign n553 = n539 ^ n537 ;
  assign n554 = n540 ^ n538 ;
  assign n555 = n553 & n554 ;
  assign n557 = n555 ^ n551 ;
  assign n546 = n535 ^ n533 ;
  assign n547 = n536 ^ n534 ;
  assign n548 = n546 & n547 ;
  assign n550 = n548 ^ n544 ;
  assign n571 = n557 ^ n550 ;
  assign n582 = n577 ^ n571 ;
  assign n583 = n582 ^ n532 ;
  assign n854 = n702 ^ n583 ;
  assign n268 = n254 ^ n252 ;
  assign n269 = n255 ^ n253 ;
  assign n270 = n268 & n269 ;
  assign n272 = n270 ^ n266 ;
  assign n261 = n250 ^ n248 ;
  assign n262 = n251 ^ n249 ;
  assign n263 = n261 & n262 ;
  assign n265 = n263 ^ n259 ;
  assign n286 = n272 ^ n265 ;
  assign n297 = n292 ^ n286 ;
  assign n298 = n297 ^ n247 ;
  assign n149 = n135 ^ n133 ;
  assign n150 = n136 ^ n134 ;
  assign n151 = n149 & n150 ;
  assign n153 = n151 ^ n147 ;
  assign n142 = n131 ^ n129 ;
  assign n143 = n132 ^ n130 ;
  assign n144 = n142 & n143 ;
  assign n146 = n144 ^ n140 ;
  assign n167 = n153 ^ n146 ;
  assign n178 = n173 ^ n167 ;
  assign n179 = n178 ^ n128 ;
  assign n450 = n298 ^ n179 ;
  assign n1329 = n854 ^ n450 ;
  assign n679 = n658 ^ n654 ;
  assign n680 = n659 ^ n655 ;
  assign n683 = n679 & n680 ;
  assign n677 = n656 ^ n652 ;
  assign n678 = n657 ^ n653 ;
  assign n682 = n677 & n678 ;
  assign n687 = n683 ^ n682 ;
  assign n691 = n689 ^ n687 ;
  assign n692 = n691 ^ n676 ;
  assign n703 = n697 ^ n692 ;
  assign n661 = n651 ^ n646 ;
  assign n704 = n703 ^ n661 ;
  assign n560 = n539 ^ n535 ;
  assign n561 = n540 ^ n536 ;
  assign n564 = n560 & n561 ;
  assign n558 = n537 ^ n533 ;
  assign n559 = n538 ^ n534 ;
  assign n563 = n558 & n559 ;
  assign n568 = n564 ^ n563 ;
  assign n572 = n570 ^ n568 ;
  assign n573 = n572 ^ n557 ;
  assign n584 = n578 ^ n573 ;
  assign n542 = n532 ^ n527 ;
  assign n585 = n584 ^ n542 ;
  assign n855 = n704 ^ n585 ;
  assign n275 = n254 ^ n250 ;
  assign n276 = n255 ^ n251 ;
  assign n279 = n275 & n276 ;
  assign n273 = n252 ^ n248 ;
  assign n274 = n253 ^ n249 ;
  assign n278 = n273 & n274 ;
  assign n283 = n279 ^ n278 ;
  assign n287 = n285 ^ n283 ;
  assign n288 = n287 ^ n272 ;
  assign n299 = n293 ^ n288 ;
  assign n257 = n247 ^ n242 ;
  assign n300 = n299 ^ n257 ;
  assign n156 = n135 ^ n131 ;
  assign n157 = n136 ^ n132 ;
  assign n160 = n156 & n157 ;
  assign n154 = n133 ^ n129 ;
  assign n155 = n134 ^ n130 ;
  assign n159 = n154 & n155 ;
  assign n164 = n160 ^ n159 ;
  assign n168 = n166 ^ n164 ;
  assign n169 = n168 ^ n153 ;
  assign n180 = n174 ^ n169 ;
  assign n138 = n128 ^ n123 ;
  assign n181 = n180 ^ n138 ;
  assign n451 = n300 ^ n181 ;
  assign n1330 = n855 ^ n451 ;
  assign n684 = n679 ^ n677 ;
  assign n685 = n680 ^ n678 ;
  assign n686 = n684 & n685 ;
  assign n688 = n686 ^ n682 ;
  assign n693 = n690 ^ n688 ;
  assign n681 = n676 ^ n675 ;
  assign n694 = n693 ^ n681 ;
  assign n705 = n698 ^ n694 ;
  assign n660 = n651 ^ n649 ;
  assign n662 = n660 ^ n647 ;
  assign n706 = n705 ^ n662 ;
  assign n565 = n560 ^ n558 ;
  assign n566 = n561 ^ n559 ;
  assign n567 = n565 & n566 ;
  assign n569 = n567 ^ n563 ;
  assign n574 = n571 ^ n569 ;
  assign n562 = n557 ^ n556 ;
  assign n575 = n574 ^ n562 ;
  assign n586 = n579 ^ n575 ;
  assign n541 = n532 ^ n530 ;
  assign n543 = n541 ^ n528 ;
  assign n587 = n586 ^ n543 ;
  assign n856 = n706 ^ n587 ;
  assign n280 = n275 ^ n273 ;
  assign n281 = n276 ^ n274 ;
  assign n282 = n280 & n281 ;
  assign n284 = n282 ^ n278 ;
  assign n289 = n286 ^ n284 ;
  assign n277 = n272 ^ n271 ;
  assign n290 = n289 ^ n277 ;
  assign n301 = n294 ^ n290 ;
  assign n256 = n247 ^ n245 ;
  assign n258 = n256 ^ n243 ;
  assign n302 = n301 ^ n258 ;
  assign n161 = n156 ^ n154 ;
  assign n162 = n157 ^ n155 ;
  assign n163 = n161 & n162 ;
  assign n165 = n163 ^ n159 ;
  assign n170 = n167 ^ n165 ;
  assign n158 = n153 ^ n152 ;
  assign n171 = n170 ^ n158 ;
  assign n182 = n175 ^ n171 ;
  assign n137 = n128 ^ n126 ;
  assign n139 = n137 ^ n124 ;
  assign n183 = n182 ^ n139 ;
  assign n452 = n302 ^ n183 ;
  assign n1331 = n856 ^ n452 ;
  assign n721 = x31 ^ x23 ;
  assign n722 = x63 ^ x55 ;
  assign n770 = n721 & n722 ;
  assign n719 = x30 ^ x22 ;
  assign n720 = x62 ^ x54 ;
  assign n769 = n719 & n720 ;
  assign n774 = n770 ^ n769 ;
  assign n717 = x29 ^ x21 ;
  assign n718 = x61 ^ x53 ;
  assign n763 = n717 & n718 ;
  assign n715 = x28 ^ x20 ;
  assign n716 = x60 ^ x52 ;
  assign n762 = n715 & n716 ;
  assign n767 = n763 ^ n762 ;
  assign n788 = n774 ^ n767 ;
  assign n713 = x27 ^ x19 ;
  assign n714 = x59 ^ x51 ;
  assign n738 = n713 & n714 ;
  assign n711 = x26 ^ x18 ;
  assign n712 = x58 ^ x50 ;
  assign n737 = n711 & n712 ;
  assign n742 = n738 ^ n737 ;
  assign n709 = x25 ^ x17 ;
  assign n710 = x57 ^ x49 ;
  assign n731 = n709 & n710 ;
  assign n707 = x24 ^ x16 ;
  assign n708 = x56 ^ x48 ;
  assign n730 = n707 & n708 ;
  assign n735 = n731 ^ n730 ;
  assign n756 = n742 ^ n735 ;
  assign n837 = n788 ^ n756 ;
  assign n857 = n849 ^ n837 ;
  assign n858 = n857 ^ n700 ;
  assign n317 = x15 ^ x7 ;
  assign n318 = x47 ^ x39 ;
  assign n366 = n317 & n318 ;
  assign n315 = x14 ^ x6 ;
  assign n316 = x46 ^ x38 ;
  assign n365 = n315 & n316 ;
  assign n370 = n366 ^ n365 ;
  assign n313 = x13 ^ x5 ;
  assign n314 = x45 ^ x37 ;
  assign n359 = n313 & n314 ;
  assign n311 = x12 ^ x4 ;
  assign n312 = x44 ^ x36 ;
  assign n358 = n311 & n312 ;
  assign n363 = n359 ^ n358 ;
  assign n384 = n370 ^ n363 ;
  assign n309 = x11 ^ x3 ;
  assign n310 = x43 ^ x35 ;
  assign n334 = n309 & n310 ;
  assign n307 = x10 ^ x2 ;
  assign n308 = x42 ^ x34 ;
  assign n333 = n307 & n308 ;
  assign n338 = n334 ^ n333 ;
  assign n305 = x9 ^ x1 ;
  assign n306 = x41 ^ x33 ;
  assign n327 = n305 & n306 ;
  assign n303 = x8 ^ x0 ;
  assign n304 = x40 ^ x32 ;
  assign n326 = n303 & n304 ;
  assign n331 = n327 ^ n326 ;
  assign n352 = n338 ^ n331 ;
  assign n433 = n384 ^ n352 ;
  assign n453 = n445 ^ n433 ;
  assign n454 = n453 ^ n296 ;
  assign n1332 = n858 ^ n454 ;
  assign n771 = n721 ^ n719 ;
  assign n772 = n722 ^ n720 ;
  assign n773 = n771 & n772 ;
  assign n775 = n773 ^ n769 ;
  assign n764 = n717 ^ n715 ;
  assign n765 = n718 ^ n716 ;
  assign n766 = n764 & n765 ;
  assign n768 = n766 ^ n762 ;
  assign n789 = n775 ^ n768 ;
  assign n739 = n713 ^ n711 ;
  assign n740 = n714 ^ n712 ;
  assign n741 = n739 & n740 ;
  assign n743 = n741 ^ n737 ;
  assign n732 = n709 ^ n707 ;
  assign n733 = n710 ^ n708 ;
  assign n734 = n732 & n733 ;
  assign n736 = n734 ^ n730 ;
  assign n757 = n743 ^ n736 ;
  assign n838 = n789 ^ n757 ;
  assign n859 = n850 ^ n838 ;
  assign n860 = n859 ^ n702 ;
  assign n367 = n317 ^ n315 ;
  assign n368 = n318 ^ n316 ;
  assign n369 = n367 & n368 ;
  assign n371 = n369 ^ n365 ;
  assign n360 = n313 ^ n311 ;
  assign n361 = n314 ^ n312 ;
  assign n362 = n360 & n361 ;
  assign n364 = n362 ^ n358 ;
  assign n385 = n371 ^ n364 ;
  assign n335 = n309 ^ n307 ;
  assign n336 = n310 ^ n308 ;
  assign n337 = n335 & n336 ;
  assign n339 = n337 ^ n333 ;
  assign n328 = n305 ^ n303 ;
  assign n329 = n306 ^ n304 ;
  assign n330 = n328 & n329 ;
  assign n332 = n330 ^ n326 ;
  assign n353 = n339 ^ n332 ;
  assign n434 = n385 ^ n353 ;
  assign n455 = n446 ^ n434 ;
  assign n456 = n455 ^ n298 ;
  assign n1333 = n860 ^ n456 ;
  assign n778 = n721 ^ n717 ;
  assign n779 = n722 ^ n718 ;
  assign n782 = n778 & n779 ;
  assign n776 = n719 ^ n715 ;
  assign n777 = n720 ^ n716 ;
  assign n781 = n776 & n777 ;
  assign n786 = n782 ^ n781 ;
  assign n790 = n788 ^ n786 ;
  assign n791 = n790 ^ n775 ;
  assign n746 = n713 ^ n709 ;
  assign n747 = n714 ^ n710 ;
  assign n750 = n746 & n747 ;
  assign n744 = n711 ^ n707 ;
  assign n745 = n712 ^ n708 ;
  assign n749 = n744 & n745 ;
  assign n754 = n750 ^ n749 ;
  assign n758 = n756 ^ n754 ;
  assign n759 = n758 ^ n743 ;
  assign n839 = n791 ^ n759 ;
  assign n861 = n851 ^ n839 ;
  assign n862 = n861 ^ n704 ;
  assign n374 = n317 ^ n313 ;
  assign n375 = n318 ^ n314 ;
  assign n378 = n374 & n375 ;
  assign n372 = n315 ^ n311 ;
  assign n373 = n316 ^ n312 ;
  assign n377 = n372 & n373 ;
  assign n382 = n378 ^ n377 ;
  assign n386 = n384 ^ n382 ;
  assign n387 = n386 ^ n371 ;
  assign n342 = n309 ^ n305 ;
  assign n343 = n310 ^ n306 ;
  assign n346 = n342 & n343 ;
  assign n340 = n307 ^ n303 ;
  assign n341 = n308 ^ n304 ;
  assign n345 = n340 & n341 ;
  assign n350 = n346 ^ n345 ;
  assign n354 = n352 ^ n350 ;
  assign n355 = n354 ^ n339 ;
  assign n435 = n387 ^ n355 ;
  assign n457 = n447 ^ n435 ;
  assign n458 = n457 ^ n300 ;
  assign n1334 = n862 ^ n458 ;
  assign n783 = n778 ^ n776 ;
  assign n784 = n779 ^ n777 ;
  assign n785 = n783 & n784 ;
  assign n787 = n785 ^ n781 ;
  assign n792 = n789 ^ n787 ;
  assign n780 = n775 ^ n774 ;
  assign n793 = n792 ^ n780 ;
  assign n751 = n746 ^ n744 ;
  assign n752 = n747 ^ n745 ;
  assign n753 = n751 & n752 ;
  assign n755 = n753 ^ n749 ;
  assign n760 = n757 ^ n755 ;
  assign n748 = n743 ^ n742 ;
  assign n761 = n760 ^ n748 ;
  assign n840 = n793 ^ n761 ;
  assign n863 = n852 ^ n840 ;
  assign n864 = n863 ^ n706 ;
  assign n379 = n374 ^ n372 ;
  assign n380 = n375 ^ n373 ;
  assign n381 = n379 & n380 ;
  assign n383 = n381 ^ n377 ;
  assign n388 = n385 ^ n383 ;
  assign n376 = n371 ^ n370 ;
  assign n389 = n388 ^ n376 ;
  assign n347 = n342 ^ n340 ;
  assign n348 = n343 ^ n341 ;
  assign n349 = n347 & n348 ;
  assign n351 = n349 ^ n345 ;
  assign n356 = n353 ^ n351 ;
  assign n344 = n339 ^ n338 ;
  assign n357 = n356 ^ n344 ;
  assign n436 = n389 ^ n357 ;
  assign n459 = n448 ^ n436 ;
  assign n460 = n459 ^ n302 ;
  assign n1335 = n864 ^ n460 ;
  assign n800 = n721 ^ n713 ;
  assign n801 = n722 ^ n714 ;
  assign n813 = n800 & n801 ;
  assign n798 = n719 ^ n711 ;
  assign n799 = n720 ^ n712 ;
  assign n812 = n798 & n799 ;
  assign n817 = n813 ^ n812 ;
  assign n796 = n717 ^ n709 ;
  assign n797 = n718 ^ n710 ;
  assign n806 = n796 & n797 ;
  assign n794 = n715 ^ n707 ;
  assign n795 = n716 ^ n708 ;
  assign n805 = n794 & n795 ;
  assign n810 = n806 ^ n805 ;
  assign n831 = n817 ^ n810 ;
  assign n841 = n837 ^ n831 ;
  assign n842 = n841 ^ n791 ;
  assign n865 = n853 ^ n842 ;
  assign n726 = n704 ^ n695 ;
  assign n866 = n865 ^ n726 ;
  assign n396 = n317 ^ n309 ;
  assign n397 = n318 ^ n310 ;
  assign n409 = n396 & n397 ;
  assign n394 = n315 ^ n307 ;
  assign n395 = n316 ^ n308 ;
  assign n408 = n394 & n395 ;
  assign n413 = n409 ^ n408 ;
  assign n392 = n313 ^ n305 ;
  assign n393 = n314 ^ n306 ;
  assign n402 = n392 & n393 ;
  assign n390 = n311 ^ n303 ;
  assign n391 = n312 ^ n304 ;
  assign n401 = n390 & n391 ;
  assign n406 = n402 ^ n401 ;
  assign n427 = n413 ^ n406 ;
  assign n437 = n433 ^ n427 ;
  assign n438 = n437 ^ n387 ;
  assign n461 = n449 ^ n438 ;
  assign n322 = n300 ^ n291 ;
  assign n462 = n461 ^ n322 ;
  assign n1336 = n866 ^ n462 ;
  assign n814 = n800 ^ n798 ;
  assign n815 = n801 ^ n799 ;
  assign n816 = n814 & n815 ;
  assign n818 = n816 ^ n812 ;
  assign n807 = n796 ^ n794 ;
  assign n808 = n797 ^ n795 ;
  assign n809 = n807 & n808 ;
  assign n811 = n809 ^ n805 ;
  assign n832 = n818 ^ n811 ;
  assign n843 = n838 ^ n832 ;
  assign n844 = n843 ^ n793 ;
  assign n867 = n854 ^ n844 ;
  assign n727 = n706 ^ n696 ;
  assign n868 = n867 ^ n727 ;
  assign n410 = n396 ^ n394 ;
  assign n411 = n397 ^ n395 ;
  assign n412 = n410 & n411 ;
  assign n414 = n412 ^ n408 ;
  assign n403 = n392 ^ n390 ;
  assign n404 = n393 ^ n391 ;
  assign n405 = n403 & n404 ;
  assign n407 = n405 ^ n401 ;
  assign n428 = n414 ^ n407 ;
  assign n439 = n434 ^ n428 ;
  assign n440 = n439 ^ n389 ;
  assign n463 = n450 ^ n440 ;
  assign n323 = n302 ^ n292 ;
  assign n464 = n463 ^ n323 ;
  assign n1337 = n868 ^ n464 ;
  assign n821 = n800 ^ n796 ;
  assign n822 = n801 ^ n797 ;
  assign n825 = n821 & n822 ;
  assign n819 = n798 ^ n794 ;
  assign n820 = n799 ^ n795 ;
  assign n824 = n819 & n820 ;
  assign n829 = n825 ^ n824 ;
  assign n833 = n831 ^ n829 ;
  assign n834 = n833 ^ n818 ;
  assign n845 = n839 ^ n834 ;
  assign n803 = n793 ^ n788 ;
  assign n846 = n845 ^ n803 ;
  assign n869 = n855 ^ n846 ;
  assign n724 = n706 ^ n700 ;
  assign n728 = n724 ^ n697 ;
  assign n870 = n869 ^ n728 ;
  assign n417 = n396 ^ n392 ;
  assign n418 = n397 ^ n393 ;
  assign n421 = n417 & n418 ;
  assign n415 = n394 ^ n390 ;
  assign n416 = n395 ^ n391 ;
  assign n420 = n415 & n416 ;
  assign n425 = n421 ^ n420 ;
  assign n429 = n427 ^ n425 ;
  assign n430 = n429 ^ n414 ;
  assign n441 = n435 ^ n430 ;
  assign n399 = n389 ^ n384 ;
  assign n442 = n441 ^ n399 ;
  assign n465 = n451 ^ n442 ;
  assign n320 = n302 ^ n296 ;
  assign n324 = n320 ^ n293 ;
  assign n466 = n465 ^ n324 ;
  assign n1338 = n870 ^ n466 ;
  assign n826 = n821 ^ n819 ;
  assign n827 = n822 ^ n820 ;
  assign n828 = n826 & n827 ;
  assign n830 = n828 ^ n824 ;
  assign n835 = n832 ^ n830 ;
  assign n823 = n818 ^ n817 ;
  assign n836 = n835 ^ n823 ;
  assign n847 = n840 ^ n836 ;
  assign n802 = n793 ^ n791 ;
  assign n804 = n802 ^ n789 ;
  assign n848 = n847 ^ n804 ;
  assign n871 = n856 ^ n848 ;
  assign n723 = n706 ^ n704 ;
  assign n725 = n723 ^ n702 ;
  assign n729 = n725 ^ n698 ;
  assign n872 = n871 ^ n729 ;
  assign n422 = n417 ^ n415 ;
  assign n423 = n418 ^ n416 ;
  assign n424 = n422 & n423 ;
  assign n426 = n424 ^ n420 ;
  assign n431 = n428 ^ n426 ;
  assign n419 = n414 ^ n413 ;
  assign n432 = n431 ^ n419 ;
  assign n443 = n436 ^ n432 ;
  assign n398 = n389 ^ n387 ;
  assign n400 = n398 ^ n385 ;
  assign n444 = n443 ^ n400 ;
  assign n467 = n452 ^ n444 ;
  assign n319 = n302 ^ n300 ;
  assign n321 = n319 ^ n298 ;
  assign n325 = n321 ^ n294 ;
  assign n468 = n467 ^ n325 ;
  assign n1339 = n872 ^ n468 ;
  assign n903 = x31 ^ x15 ;
  assign n904 = x63 ^ x47 ;
  assign n1079 = n903 & n904 ;
  assign n901 = x30 ^ x14 ;
  assign n902 = x62 ^ x46 ;
  assign n1078 = n901 & n902 ;
  assign n1083 = n1079 ^ n1078 ;
  assign n899 = x29 ^ x13 ;
  assign n900 = x61 ^ x45 ;
  assign n1072 = n899 & n900 ;
  assign n897 = x28 ^ x12 ;
  assign n898 = x60 ^ x44 ;
  assign n1071 = n897 & n898 ;
  assign n1076 = n1072 ^ n1071 ;
  assign n1097 = n1083 ^ n1076 ;
  assign n895 = x27 ^ x11 ;
  assign n896 = x59 ^ x43 ;
  assign n1047 = n895 & n896 ;
  assign n893 = x26 ^ x10 ;
  assign n894 = x58 ^ x42 ;
  assign n1046 = n893 & n894 ;
  assign n1051 = n1047 ^ n1046 ;
  assign n891 = x25 ^ x9 ;
  assign n892 = x57 ^ x41 ;
  assign n1040 = n891 & n892 ;
  assign n889 = x24 ^ x8 ;
  assign n890 = x56 ^ x40 ;
  assign n1039 = n889 & n890 ;
  assign n1044 = n1040 ^ n1039 ;
  assign n1065 = n1051 ^ n1044 ;
  assign n1146 = n1097 ^ n1065 ;
  assign n887 = x23 ^ x7 ;
  assign n888 = x55 ^ x39 ;
  assign n960 = n887 & n888 ;
  assign n885 = x22 ^ x6 ;
  assign n886 = x54 ^ x38 ;
  assign n959 = n885 & n886 ;
  assign n964 = n960 ^ n959 ;
  assign n883 = x21 ^ x5 ;
  assign n884 = x53 ^ x37 ;
  assign n953 = n883 & n884 ;
  assign n881 = x20 ^ x4 ;
  assign n882 = x52 ^ x36 ;
  assign n952 = n881 & n882 ;
  assign n957 = n953 ^ n952 ;
  assign n978 = n964 ^ n957 ;
  assign n879 = x19 ^ x3 ;
  assign n880 = x51 ^ x35 ;
  assign n928 = n879 & n880 ;
  assign n877 = x18 ^ x2 ;
  assign n878 = x50 ^ x34 ;
  assign n927 = n877 & n878 ;
  assign n932 = n928 ^ n927 ;
  assign n875 = x17 ^ x1 ;
  assign n876 = x49 ^ x33 ;
  assign n921 = n875 & n876 ;
  assign n873 = x16 ^ x0 ;
  assign n874 = x48 ^ x32 ;
  assign n920 = n873 & n874 ;
  assign n925 = n921 ^ n920 ;
  assign n946 = n932 ^ n925 ;
  assign n1027 = n978 ^ n946 ;
  assign n1300 = n1146 ^ n1027 ;
  assign n1340 = n1324 ^ n1300 ;
  assign n1341 = n1340 ^ n858 ;
  assign n1080 = n903 ^ n901 ;
  assign n1081 = n904 ^ n902 ;
  assign n1082 = n1080 & n1081 ;
  assign n1084 = n1082 ^ n1078 ;
  assign n1073 = n899 ^ n897 ;
  assign n1074 = n900 ^ n898 ;
  assign n1075 = n1073 & n1074 ;
  assign n1077 = n1075 ^ n1071 ;
  assign n1098 = n1084 ^ n1077 ;
  assign n1048 = n895 ^ n893 ;
  assign n1049 = n896 ^ n894 ;
  assign n1050 = n1048 & n1049 ;
  assign n1052 = n1050 ^ n1046 ;
  assign n1041 = n891 ^ n889 ;
  assign n1042 = n892 ^ n890 ;
  assign n1043 = n1041 & n1042 ;
  assign n1045 = n1043 ^ n1039 ;
  assign n1066 = n1052 ^ n1045 ;
  assign n1147 = n1098 ^ n1066 ;
  assign n961 = n887 ^ n885 ;
  assign n962 = n888 ^ n886 ;
  assign n963 = n961 & n962 ;
  assign n965 = n963 ^ n959 ;
  assign n954 = n883 ^ n881 ;
  assign n955 = n884 ^ n882 ;
  assign n956 = n954 & n955 ;
  assign n958 = n956 ^ n952 ;
  assign n979 = n965 ^ n958 ;
  assign n929 = n879 ^ n877 ;
  assign n930 = n880 ^ n878 ;
  assign n931 = n929 & n930 ;
  assign n933 = n931 ^ n927 ;
  assign n922 = n875 ^ n873 ;
  assign n923 = n876 ^ n874 ;
  assign n924 = n922 & n923 ;
  assign n926 = n924 ^ n920 ;
  assign n947 = n933 ^ n926 ;
  assign n1028 = n979 ^ n947 ;
  assign n1301 = n1147 ^ n1028 ;
  assign n1342 = n1325 ^ n1301 ;
  assign n1343 = n1342 ^ n860 ;
  assign n1087 = n903 ^ n899 ;
  assign n1088 = n904 ^ n900 ;
  assign n1091 = n1087 & n1088 ;
  assign n1085 = n901 ^ n897 ;
  assign n1086 = n902 ^ n898 ;
  assign n1090 = n1085 & n1086 ;
  assign n1095 = n1091 ^ n1090 ;
  assign n1099 = n1097 ^ n1095 ;
  assign n1100 = n1099 ^ n1084 ;
  assign n1055 = n895 ^ n891 ;
  assign n1056 = n896 ^ n892 ;
  assign n1059 = n1055 & n1056 ;
  assign n1053 = n893 ^ n889 ;
  assign n1054 = n894 ^ n890 ;
  assign n1058 = n1053 & n1054 ;
  assign n1063 = n1059 ^ n1058 ;
  assign n1067 = n1065 ^ n1063 ;
  assign n1068 = n1067 ^ n1052 ;
  assign n1148 = n1100 ^ n1068 ;
  assign n968 = n887 ^ n883 ;
  assign n969 = n888 ^ n884 ;
  assign n972 = n968 & n969 ;
  assign n966 = n885 ^ n881 ;
  assign n967 = n886 ^ n882 ;
  assign n971 = n966 & n967 ;
  assign n976 = n972 ^ n971 ;
  assign n980 = n978 ^ n976 ;
  assign n981 = n980 ^ n965 ;
  assign n936 = n879 ^ n875 ;
  assign n937 = n880 ^ n876 ;
  assign n940 = n936 & n937 ;
  assign n934 = n877 ^ n873 ;
  assign n935 = n878 ^ n874 ;
  assign n939 = n934 & n935 ;
  assign n944 = n940 ^ n939 ;
  assign n948 = n946 ^ n944 ;
  assign n949 = n948 ^ n933 ;
  assign n1029 = n981 ^ n949 ;
  assign n1302 = n1148 ^ n1029 ;
  assign n1344 = n1326 ^ n1302 ;
  assign n1345 = n1344 ^ n862 ;
  assign n1092 = n1087 ^ n1085 ;
  assign n1093 = n1088 ^ n1086 ;
  assign n1094 = n1092 & n1093 ;
  assign n1096 = n1094 ^ n1090 ;
  assign n1101 = n1098 ^ n1096 ;
  assign n1089 = n1084 ^ n1083 ;
  assign n1102 = n1101 ^ n1089 ;
  assign n1060 = n1055 ^ n1053 ;
  assign n1061 = n1056 ^ n1054 ;
  assign n1062 = n1060 & n1061 ;
  assign n1064 = n1062 ^ n1058 ;
  assign n1069 = n1066 ^ n1064 ;
  assign n1057 = n1052 ^ n1051 ;
  assign n1070 = n1069 ^ n1057 ;
  assign n1149 = n1102 ^ n1070 ;
  assign n973 = n968 ^ n966 ;
  assign n974 = n969 ^ n967 ;
  assign n975 = n973 & n974 ;
  assign n977 = n975 ^ n971 ;
  assign n982 = n979 ^ n977 ;
  assign n970 = n965 ^ n964 ;
  assign n983 = n982 ^ n970 ;
  assign n941 = n936 ^ n934 ;
  assign n942 = n937 ^ n935 ;
  assign n943 = n941 & n942 ;
  assign n945 = n943 ^ n939 ;
  assign n950 = n947 ^ n945 ;
  assign n938 = n933 ^ n932 ;
  assign n951 = n950 ^ n938 ;
  assign n1030 = n983 ^ n951 ;
  assign n1303 = n1149 ^ n1030 ;
  assign n1346 = n1327 ^ n1303 ;
  assign n1347 = n1346 ^ n864 ;
  assign n1109 = n903 ^ n895 ;
  assign n1110 = n904 ^ n896 ;
  assign n1122 = n1109 & n1110 ;
  assign n1107 = n901 ^ n893 ;
  assign n1108 = n902 ^ n894 ;
  assign n1121 = n1107 & n1108 ;
  assign n1126 = n1122 ^ n1121 ;
  assign n1105 = n899 ^ n891 ;
  assign n1106 = n900 ^ n892 ;
  assign n1115 = n1105 & n1106 ;
  assign n1103 = n897 ^ n889 ;
  assign n1104 = n898 ^ n890 ;
  assign n1114 = n1103 & n1104 ;
  assign n1119 = n1115 ^ n1114 ;
  assign n1140 = n1126 ^ n1119 ;
  assign n1150 = n1146 ^ n1140 ;
  assign n1151 = n1150 ^ n1100 ;
  assign n990 = n887 ^ n879 ;
  assign n991 = n888 ^ n880 ;
  assign n1003 = n990 & n991 ;
  assign n988 = n885 ^ n877 ;
  assign n989 = n886 ^ n878 ;
  assign n1002 = n988 & n989 ;
  assign n1007 = n1003 ^ n1002 ;
  assign n986 = n883 ^ n875 ;
  assign n987 = n884 ^ n876 ;
  assign n996 = n986 & n987 ;
  assign n984 = n881 ^ n873 ;
  assign n985 = n882 ^ n874 ;
  assign n995 = n984 & n985 ;
  assign n1000 = n996 ^ n995 ;
  assign n1021 = n1007 ^ n1000 ;
  assign n1031 = n1027 ^ n1021 ;
  assign n1032 = n1031 ^ n981 ;
  assign n1304 = n1151 ^ n1032 ;
  assign n1348 = n1328 ^ n1304 ;
  assign n1349 = n1348 ^ n866 ;
  assign n1123 = n1109 ^ n1107 ;
  assign n1124 = n1110 ^ n1108 ;
  assign n1125 = n1123 & n1124 ;
  assign n1127 = n1125 ^ n1121 ;
  assign n1116 = n1105 ^ n1103 ;
  assign n1117 = n1106 ^ n1104 ;
  assign n1118 = n1116 & n1117 ;
  assign n1120 = n1118 ^ n1114 ;
  assign n1141 = n1127 ^ n1120 ;
  assign n1152 = n1147 ^ n1141 ;
  assign n1153 = n1152 ^ n1102 ;
  assign n1004 = n990 ^ n988 ;
  assign n1005 = n991 ^ n989 ;
  assign n1006 = n1004 & n1005 ;
  assign n1008 = n1006 ^ n1002 ;
  assign n997 = n986 ^ n984 ;
  assign n998 = n987 ^ n985 ;
  assign n999 = n997 & n998 ;
  assign n1001 = n999 ^ n995 ;
  assign n1022 = n1008 ^ n1001 ;
  assign n1033 = n1028 ^ n1022 ;
  assign n1034 = n1033 ^ n983 ;
  assign n1305 = n1153 ^ n1034 ;
  assign n1350 = n1329 ^ n1305 ;
  assign n1351 = n1350 ^ n868 ;
  assign n1130 = n1109 ^ n1105 ;
  assign n1131 = n1110 ^ n1106 ;
  assign n1134 = n1130 & n1131 ;
  assign n1128 = n1107 ^ n1103 ;
  assign n1129 = n1108 ^ n1104 ;
  assign n1133 = n1128 & n1129 ;
  assign n1138 = n1134 ^ n1133 ;
  assign n1142 = n1140 ^ n1138 ;
  assign n1143 = n1142 ^ n1127 ;
  assign n1154 = n1148 ^ n1143 ;
  assign n1112 = n1102 ^ n1097 ;
  assign n1155 = n1154 ^ n1112 ;
  assign n1011 = n990 ^ n986 ;
  assign n1012 = n991 ^ n987 ;
  assign n1015 = n1011 & n1012 ;
  assign n1009 = n988 ^ n984 ;
  assign n1010 = n989 ^ n985 ;
  assign n1014 = n1009 & n1010 ;
  assign n1019 = n1015 ^ n1014 ;
  assign n1023 = n1021 ^ n1019 ;
  assign n1024 = n1023 ^ n1008 ;
  assign n1035 = n1029 ^ n1024 ;
  assign n993 = n983 ^ n978 ;
  assign n1036 = n1035 ^ n993 ;
  assign n1306 = n1155 ^ n1036 ;
  assign n1352 = n1330 ^ n1306 ;
  assign n1353 = n1352 ^ n870 ;
  assign n1135 = n1130 ^ n1128 ;
  assign n1136 = n1131 ^ n1129 ;
  assign n1137 = n1135 & n1136 ;
  assign n1139 = n1137 ^ n1133 ;
  assign n1144 = n1141 ^ n1139 ;
  assign n1132 = n1127 ^ n1126 ;
  assign n1145 = n1144 ^ n1132 ;
  assign n1156 = n1149 ^ n1145 ;
  assign n1111 = n1102 ^ n1100 ;
  assign n1113 = n1111 ^ n1098 ;
  assign n1157 = n1156 ^ n1113 ;
  assign n1016 = n1011 ^ n1009 ;
  assign n1017 = n1012 ^ n1010 ;
  assign n1018 = n1016 & n1017 ;
  assign n1020 = n1018 ^ n1014 ;
  assign n1025 = n1022 ^ n1020 ;
  assign n1013 = n1008 ^ n1007 ;
  assign n1026 = n1025 ^ n1013 ;
  assign n1037 = n1030 ^ n1026 ;
  assign n992 = n983 ^ n981 ;
  assign n994 = n992 ^ n979 ;
  assign n1038 = n1037 ^ n994 ;
  assign n1307 = n1157 ^ n1038 ;
  assign n1354 = n1331 ^ n1307 ;
  assign n1355 = n1354 ^ n872 ;
  assign n1172 = n903 ^ n887 ;
  assign n1173 = n904 ^ n888 ;
  assign n1221 = n1172 & n1173 ;
  assign n1170 = n901 ^ n885 ;
  assign n1171 = n902 ^ n886 ;
  assign n1220 = n1170 & n1171 ;
  assign n1225 = n1221 ^ n1220 ;
  assign n1168 = n899 ^ n883 ;
  assign n1169 = n900 ^ n884 ;
  assign n1214 = n1168 & n1169 ;
  assign n1166 = n897 ^ n881 ;
  assign n1167 = n898 ^ n882 ;
  assign n1213 = n1166 & n1167 ;
  assign n1218 = n1214 ^ n1213 ;
  assign n1239 = n1225 ^ n1218 ;
  assign n1164 = n895 ^ n879 ;
  assign n1165 = n896 ^ n880 ;
  assign n1189 = n1164 & n1165 ;
  assign n1162 = n893 ^ n877 ;
  assign n1163 = n894 ^ n878 ;
  assign n1188 = n1162 & n1163 ;
  assign n1193 = n1189 ^ n1188 ;
  assign n1160 = n891 ^ n875 ;
  assign n1161 = n892 ^ n876 ;
  assign n1182 = n1160 & n1161 ;
  assign n1158 = n889 ^ n873 ;
  assign n1159 = n890 ^ n874 ;
  assign n1181 = n1158 & n1159 ;
  assign n1186 = n1182 ^ n1181 ;
  assign n1207 = n1193 ^ n1186 ;
  assign n1288 = n1239 ^ n1207 ;
  assign n1308 = n1300 ^ n1288 ;
  assign n1309 = n1308 ^ n1151 ;
  assign n1356 = n1332 ^ n1309 ;
  assign n912 = n866 ^ n849 ;
  assign n1357 = n1356 ^ n912 ;
  assign n1222 = n1172 ^ n1170 ;
  assign n1223 = n1173 ^ n1171 ;
  assign n1224 = n1222 & n1223 ;
  assign n1226 = n1224 ^ n1220 ;
  assign n1215 = n1168 ^ n1166 ;
  assign n1216 = n1169 ^ n1167 ;
  assign n1217 = n1215 & n1216 ;
  assign n1219 = n1217 ^ n1213 ;
  assign n1240 = n1226 ^ n1219 ;
  assign n1190 = n1164 ^ n1162 ;
  assign n1191 = n1165 ^ n1163 ;
  assign n1192 = n1190 & n1191 ;
  assign n1194 = n1192 ^ n1188 ;
  assign n1183 = n1160 ^ n1158 ;
  assign n1184 = n1161 ^ n1159 ;
  assign n1185 = n1183 & n1184 ;
  assign n1187 = n1185 ^ n1181 ;
  assign n1208 = n1194 ^ n1187 ;
  assign n1289 = n1240 ^ n1208 ;
  assign n1310 = n1301 ^ n1289 ;
  assign n1311 = n1310 ^ n1153 ;
  assign n1358 = n1333 ^ n1311 ;
  assign n913 = n868 ^ n850 ;
  assign n1359 = n1358 ^ n913 ;
  assign n1229 = n1172 ^ n1168 ;
  assign n1230 = n1173 ^ n1169 ;
  assign n1233 = n1229 & n1230 ;
  assign n1227 = n1170 ^ n1166 ;
  assign n1228 = n1171 ^ n1167 ;
  assign n1232 = n1227 & n1228 ;
  assign n1237 = n1233 ^ n1232 ;
  assign n1241 = n1239 ^ n1237 ;
  assign n1242 = n1241 ^ n1226 ;
  assign n1197 = n1164 ^ n1160 ;
  assign n1198 = n1165 ^ n1161 ;
  assign n1201 = n1197 & n1198 ;
  assign n1195 = n1162 ^ n1158 ;
  assign n1196 = n1163 ^ n1159 ;
  assign n1200 = n1195 & n1196 ;
  assign n1205 = n1201 ^ n1200 ;
  assign n1209 = n1207 ^ n1205 ;
  assign n1210 = n1209 ^ n1194 ;
  assign n1290 = n1242 ^ n1210 ;
  assign n1312 = n1302 ^ n1290 ;
  assign n1313 = n1312 ^ n1155 ;
  assign n1360 = n1334 ^ n1313 ;
  assign n914 = n870 ^ n851 ;
  assign n1361 = n1360 ^ n914 ;
  assign n1234 = n1229 ^ n1227 ;
  assign n1235 = n1230 ^ n1228 ;
  assign n1236 = n1234 & n1235 ;
  assign n1238 = n1236 ^ n1232 ;
  assign n1243 = n1240 ^ n1238 ;
  assign n1231 = n1226 ^ n1225 ;
  assign n1244 = n1243 ^ n1231 ;
  assign n1202 = n1197 ^ n1195 ;
  assign n1203 = n1198 ^ n1196 ;
  assign n1204 = n1202 & n1203 ;
  assign n1206 = n1204 ^ n1200 ;
  assign n1211 = n1208 ^ n1206 ;
  assign n1199 = n1194 ^ n1193 ;
  assign n1212 = n1211 ^ n1199 ;
  assign n1291 = n1244 ^ n1212 ;
  assign n1314 = n1303 ^ n1291 ;
  assign n1315 = n1314 ^ n1157 ;
  assign n1362 = n1335 ^ n1315 ;
  assign n915 = n872 ^ n852 ;
  assign n1363 = n1362 ^ n915 ;
  assign n1251 = n1172 ^ n1164 ;
  assign n1252 = n1173 ^ n1165 ;
  assign n1264 = n1251 & n1252 ;
  assign n1249 = n1170 ^ n1162 ;
  assign n1250 = n1171 ^ n1163 ;
  assign n1263 = n1249 & n1250 ;
  assign n1268 = n1264 ^ n1263 ;
  assign n1247 = n1168 ^ n1160 ;
  assign n1248 = n1169 ^ n1161 ;
  assign n1257 = n1247 & n1248 ;
  assign n1245 = n1166 ^ n1158 ;
  assign n1246 = n1167 ^ n1159 ;
  assign n1256 = n1245 & n1246 ;
  assign n1261 = n1257 ^ n1256 ;
  assign n1282 = n1268 ^ n1261 ;
  assign n1292 = n1288 ^ n1282 ;
  assign n1293 = n1292 ^ n1242 ;
  assign n1316 = n1304 ^ n1293 ;
  assign n1177 = n1155 ^ n1146 ;
  assign n1317 = n1316 ^ n1177 ;
  assign n1364 = n1336 ^ n1317 ;
  assign n908 = n870 ^ n858 ;
  assign n916 = n908 ^ n853 ;
  assign n1365 = n1364 ^ n916 ;
  assign n1265 = n1251 ^ n1249 ;
  assign n1266 = n1252 ^ n1250 ;
  assign n1267 = n1265 & n1266 ;
  assign n1269 = n1267 ^ n1263 ;
  assign n1258 = n1247 ^ n1245 ;
  assign n1259 = n1248 ^ n1246 ;
  assign n1260 = n1258 & n1259 ;
  assign n1262 = n1260 ^ n1256 ;
  assign n1283 = n1269 ^ n1262 ;
  assign n1294 = n1289 ^ n1283 ;
  assign n1295 = n1294 ^ n1244 ;
  assign n1318 = n1305 ^ n1295 ;
  assign n1178 = n1157 ^ n1147 ;
  assign n1319 = n1318 ^ n1178 ;
  assign n1366 = n1337 ^ n1319 ;
  assign n909 = n872 ^ n860 ;
  assign n917 = n909 ^ n854 ;
  assign n1367 = n1366 ^ n917 ;
  assign n1272 = n1251 ^ n1247 ;
  assign n1273 = n1252 ^ n1248 ;
  assign n1276 = n1272 & n1273 ;
  assign n1270 = n1249 ^ n1245 ;
  assign n1271 = n1250 ^ n1246 ;
  assign n1275 = n1270 & n1271 ;
  assign n1280 = n1276 ^ n1275 ;
  assign n1284 = n1282 ^ n1280 ;
  assign n1285 = n1284 ^ n1269 ;
  assign n1296 = n1290 ^ n1285 ;
  assign n1254 = n1244 ^ n1239 ;
  assign n1297 = n1296 ^ n1254 ;
  assign n1320 = n1306 ^ n1297 ;
  assign n1175 = n1157 ^ n1151 ;
  assign n1179 = n1175 ^ n1148 ;
  assign n1321 = n1320 ^ n1179 ;
  assign n1368 = n1338 ^ n1321 ;
  assign n906 = n872 ^ n866 ;
  assign n910 = n906 ^ n862 ;
  assign n918 = n910 ^ n855 ;
  assign n1369 = n1368 ^ n918 ;
  assign n1277 = n1272 ^ n1270 ;
  assign n1278 = n1273 ^ n1271 ;
  assign n1279 = n1277 & n1278 ;
  assign n1281 = n1279 ^ n1275 ;
  assign n1286 = n1283 ^ n1281 ;
  assign n1274 = n1269 ^ n1268 ;
  assign n1287 = n1286 ^ n1274 ;
  assign n1298 = n1291 ^ n1287 ;
  assign n1253 = n1244 ^ n1242 ;
  assign n1255 = n1253 ^ n1240 ;
  assign n1299 = n1298 ^ n1255 ;
  assign n1322 = n1307 ^ n1299 ;
  assign n1174 = n1157 ^ n1155 ;
  assign n1176 = n1174 ^ n1153 ;
  assign n1180 = n1176 ^ n1149 ;
  assign n1323 = n1322 ^ n1180 ;
  assign n1370 = n1339 ^ n1323 ;
  assign n905 = n872 ^ n870 ;
  assign n907 = n905 ^ n868 ;
  assign n911 = n907 ^ n864 ;
  assign n919 = n911 ^ n856 ;
  assign n1371 = n1370 ^ n919 ;
  assign y0 = n1324 ;
  assign y1 = n1325 ;
  assign y2 = n1326 ;
  assign y3 = n1327 ;
  assign y4 = n1328 ;
  assign y5 = n1329 ;
  assign y6 = n1330 ;
  assign y7 = n1331 ;
  assign y8 = n1332 ;
  assign y9 = n1333 ;
  assign y10 = n1334 ;
  assign y11 = n1335 ;
  assign y12 = n1336 ;
  assign y13 = n1337 ;
  assign y14 = n1338 ;
  assign y15 = n1339 ;
  assign y16 = n1341 ;
  assign y17 = n1343 ;
  assign y18 = n1345 ;
  assign y19 = n1347 ;
  assign y20 = n1349 ;
  assign y21 = n1351 ;
  assign y22 = n1353 ;
  assign y23 = n1355 ;
  assign y24 = n1357 ;
  assign y25 = n1359 ;
  assign y26 = n1361 ;
  assign y27 = n1363 ;
  assign y28 = n1365 ;
  assign y29 = n1367 ;
  assign y30 = n1369 ;
  assign y31 = n1371 ;
endmodule
