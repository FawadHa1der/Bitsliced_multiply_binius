module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 ;
  assign n192 = x15 & x31 ;
  assign n191 = x14 & x30 ;
  assign n196 = n192 ^ n191 ;
  assign n185 = x13 & x29 ;
  assign n184 = x12 & x28 ;
  assign n189 = n185 ^ n184 ;
  assign n210 = n196 ^ n189 ;
  assign n160 = x11 & x27 ;
  assign n159 = x10 & x26 ;
  assign n164 = n160 ^ n159 ;
  assign n153 = x9 & x25 ;
  assign n152 = x8 & x24 ;
  assign n157 = n153 ^ n152 ;
  assign n178 = n164 ^ n157 ;
  assign n259 = n210 ^ n178 ;
  assign n73 = x7 & x23 ;
  assign n72 = x6 & x22 ;
  assign n77 = n73 ^ n72 ;
  assign n66 = x5 & x21 ;
  assign n65 = x4 & x20 ;
  assign n70 = n66 ^ n65 ;
  assign n91 = n77 ^ n70 ;
  assign n41 = x3 & x19 ;
  assign n40 = x2 & x18 ;
  assign n45 = n41 ^ n40 ;
  assign n34 = x1 & x17 ;
  assign n33 = x0 & x16 ;
  assign n38 = n34 ^ n33 ;
  assign n59 = n45 ^ n38 ;
  assign n140 = n91 ^ n59 ;
  assign n413 = n259 ^ n140 ;
  assign n193 = x15 ^ x14 ;
  assign n194 = x31 ^ x30 ;
  assign n195 = n193 & n194 ;
  assign n197 = n195 ^ n191 ;
  assign n186 = x13 ^ x12 ;
  assign n187 = x29 ^ x28 ;
  assign n188 = n186 & n187 ;
  assign n190 = n188 ^ n184 ;
  assign n211 = n197 ^ n190 ;
  assign n161 = x11 ^ x10 ;
  assign n162 = x27 ^ x26 ;
  assign n163 = n161 & n162 ;
  assign n165 = n163 ^ n159 ;
  assign n154 = x9 ^ x8 ;
  assign n155 = x25 ^ x24 ;
  assign n156 = n154 & n155 ;
  assign n158 = n156 ^ n152 ;
  assign n179 = n165 ^ n158 ;
  assign n260 = n211 ^ n179 ;
  assign n74 = x7 ^ x6 ;
  assign n75 = x23 ^ x22 ;
  assign n76 = n74 & n75 ;
  assign n78 = n76 ^ n72 ;
  assign n67 = x5 ^ x4 ;
  assign n68 = x21 ^ x20 ;
  assign n69 = n67 & n68 ;
  assign n71 = n69 ^ n65 ;
  assign n92 = n78 ^ n71 ;
  assign n42 = x3 ^ x2 ;
  assign n43 = x19 ^ x18 ;
  assign n44 = n42 & n43 ;
  assign n46 = n44 ^ n40 ;
  assign n35 = x1 ^ x0 ;
  assign n36 = x17 ^ x16 ;
  assign n37 = n35 & n36 ;
  assign n39 = n37 ^ n33 ;
  assign n60 = n46 ^ n39 ;
  assign n141 = n92 ^ n60 ;
  assign n414 = n260 ^ n141 ;
  assign n200 = x15 ^ x13 ;
  assign n201 = x31 ^ x29 ;
  assign n204 = n200 & n201 ;
  assign n198 = x14 ^ x12 ;
  assign n199 = x30 ^ x28 ;
  assign n203 = n198 & n199 ;
  assign n208 = n204 ^ n203 ;
  assign n212 = n210 ^ n208 ;
  assign n213 = n212 ^ n197 ;
  assign n168 = x11 ^ x9 ;
  assign n169 = x27 ^ x25 ;
  assign n172 = n168 & n169 ;
  assign n166 = x10 ^ x8 ;
  assign n167 = x26 ^ x24 ;
  assign n171 = n166 & n167 ;
  assign n176 = n172 ^ n171 ;
  assign n180 = n178 ^ n176 ;
  assign n181 = n180 ^ n165 ;
  assign n261 = n213 ^ n181 ;
  assign n81 = x7 ^ x5 ;
  assign n82 = x23 ^ x21 ;
  assign n85 = n81 & n82 ;
  assign n79 = x6 ^ x4 ;
  assign n80 = x22 ^ x20 ;
  assign n84 = n79 & n80 ;
  assign n89 = n85 ^ n84 ;
  assign n93 = n91 ^ n89 ;
  assign n94 = n93 ^ n78 ;
  assign n49 = x3 ^ x1 ;
  assign n50 = x19 ^ x17 ;
  assign n53 = n49 & n50 ;
  assign n47 = x2 ^ x0 ;
  assign n48 = x18 ^ x16 ;
  assign n52 = n47 & n48 ;
  assign n57 = n53 ^ n52 ;
  assign n61 = n59 ^ n57 ;
  assign n62 = n61 ^ n46 ;
  assign n142 = n94 ^ n62 ;
  assign n415 = n261 ^ n142 ;
  assign n205 = n200 ^ n198 ;
  assign n206 = n201 ^ n199 ;
  assign n207 = n205 & n206 ;
  assign n209 = n207 ^ n203 ;
  assign n214 = n211 ^ n209 ;
  assign n202 = n197 ^ n196 ;
  assign n215 = n214 ^ n202 ;
  assign n173 = n168 ^ n166 ;
  assign n174 = n169 ^ n167 ;
  assign n175 = n173 & n174 ;
  assign n177 = n175 ^ n171 ;
  assign n182 = n179 ^ n177 ;
  assign n170 = n165 ^ n164 ;
  assign n183 = n182 ^ n170 ;
  assign n262 = n215 ^ n183 ;
  assign n86 = n81 ^ n79 ;
  assign n87 = n82 ^ n80 ;
  assign n88 = n86 & n87 ;
  assign n90 = n88 ^ n84 ;
  assign n95 = n92 ^ n90 ;
  assign n83 = n78 ^ n77 ;
  assign n96 = n95 ^ n83 ;
  assign n54 = n49 ^ n47 ;
  assign n55 = n50 ^ n48 ;
  assign n56 = n54 & n55 ;
  assign n58 = n56 ^ n52 ;
  assign n63 = n60 ^ n58 ;
  assign n51 = n46 ^ n45 ;
  assign n64 = n63 ^ n51 ;
  assign n143 = n96 ^ n64 ;
  assign n416 = n262 ^ n143 ;
  assign n222 = x15 ^ x11 ;
  assign n223 = x31 ^ x27 ;
  assign n235 = n222 & n223 ;
  assign n220 = x14 ^ x10 ;
  assign n221 = x30 ^ x26 ;
  assign n234 = n220 & n221 ;
  assign n239 = n235 ^ n234 ;
  assign n218 = x13 ^ x9 ;
  assign n219 = x29 ^ x25 ;
  assign n228 = n218 & n219 ;
  assign n216 = x12 ^ x8 ;
  assign n217 = x28 ^ x24 ;
  assign n227 = n216 & n217 ;
  assign n232 = n228 ^ n227 ;
  assign n253 = n239 ^ n232 ;
  assign n263 = n259 ^ n253 ;
  assign n264 = n263 ^ n213 ;
  assign n103 = x7 ^ x3 ;
  assign n104 = x23 ^ x19 ;
  assign n116 = n103 & n104 ;
  assign n101 = x6 ^ x2 ;
  assign n102 = x22 ^ x18 ;
  assign n115 = n101 & n102 ;
  assign n120 = n116 ^ n115 ;
  assign n99 = x5 ^ x1 ;
  assign n100 = x21 ^ x17 ;
  assign n109 = n99 & n100 ;
  assign n97 = x4 ^ x0 ;
  assign n98 = x20 ^ x16 ;
  assign n108 = n97 & n98 ;
  assign n113 = n109 ^ n108 ;
  assign n134 = n120 ^ n113 ;
  assign n144 = n140 ^ n134 ;
  assign n145 = n144 ^ n94 ;
  assign n417 = n264 ^ n145 ;
  assign n236 = n222 ^ n220 ;
  assign n237 = n223 ^ n221 ;
  assign n238 = n236 & n237 ;
  assign n240 = n238 ^ n234 ;
  assign n229 = n218 ^ n216 ;
  assign n230 = n219 ^ n217 ;
  assign n231 = n229 & n230 ;
  assign n233 = n231 ^ n227 ;
  assign n254 = n240 ^ n233 ;
  assign n265 = n260 ^ n254 ;
  assign n266 = n265 ^ n215 ;
  assign n117 = n103 ^ n101 ;
  assign n118 = n104 ^ n102 ;
  assign n119 = n117 & n118 ;
  assign n121 = n119 ^ n115 ;
  assign n110 = n99 ^ n97 ;
  assign n111 = n100 ^ n98 ;
  assign n112 = n110 & n111 ;
  assign n114 = n112 ^ n108 ;
  assign n135 = n121 ^ n114 ;
  assign n146 = n141 ^ n135 ;
  assign n147 = n146 ^ n96 ;
  assign n418 = n266 ^ n147 ;
  assign n243 = n222 ^ n218 ;
  assign n244 = n223 ^ n219 ;
  assign n247 = n243 & n244 ;
  assign n241 = n220 ^ n216 ;
  assign n242 = n221 ^ n217 ;
  assign n246 = n241 & n242 ;
  assign n251 = n247 ^ n246 ;
  assign n255 = n253 ^ n251 ;
  assign n256 = n255 ^ n240 ;
  assign n267 = n261 ^ n256 ;
  assign n225 = n215 ^ n210 ;
  assign n268 = n267 ^ n225 ;
  assign n124 = n103 ^ n99 ;
  assign n125 = n104 ^ n100 ;
  assign n128 = n124 & n125 ;
  assign n122 = n101 ^ n97 ;
  assign n123 = n102 ^ n98 ;
  assign n127 = n122 & n123 ;
  assign n132 = n128 ^ n127 ;
  assign n136 = n134 ^ n132 ;
  assign n137 = n136 ^ n121 ;
  assign n148 = n142 ^ n137 ;
  assign n106 = n96 ^ n91 ;
  assign n149 = n148 ^ n106 ;
  assign n419 = n268 ^ n149 ;
  assign n248 = n243 ^ n241 ;
  assign n249 = n244 ^ n242 ;
  assign n250 = n248 & n249 ;
  assign n252 = n250 ^ n246 ;
  assign n257 = n254 ^ n252 ;
  assign n245 = n240 ^ n239 ;
  assign n258 = n257 ^ n245 ;
  assign n269 = n262 ^ n258 ;
  assign n224 = n215 ^ n213 ;
  assign n226 = n224 ^ n211 ;
  assign n270 = n269 ^ n226 ;
  assign n129 = n124 ^ n122 ;
  assign n130 = n125 ^ n123 ;
  assign n131 = n129 & n130 ;
  assign n133 = n131 ^ n127 ;
  assign n138 = n135 ^ n133 ;
  assign n126 = n121 ^ n120 ;
  assign n139 = n138 ^ n126 ;
  assign n150 = n143 ^ n139 ;
  assign n105 = n96 ^ n94 ;
  assign n107 = n105 ^ n92 ;
  assign n151 = n150 ^ n107 ;
  assign n420 = n270 ^ n151 ;
  assign n285 = x15 ^ x7 ;
  assign n286 = x31 ^ x23 ;
  assign n334 = n285 & n286 ;
  assign n283 = x14 ^ x6 ;
  assign n284 = x30 ^ x22 ;
  assign n333 = n283 & n284 ;
  assign n338 = n334 ^ n333 ;
  assign n281 = x13 ^ x5 ;
  assign n282 = x29 ^ x21 ;
  assign n327 = n281 & n282 ;
  assign n279 = x12 ^ x4 ;
  assign n280 = x28 ^ x20 ;
  assign n326 = n279 & n280 ;
  assign n331 = n327 ^ n326 ;
  assign n352 = n338 ^ n331 ;
  assign n277 = x11 ^ x3 ;
  assign n278 = x27 ^ x19 ;
  assign n302 = n277 & n278 ;
  assign n275 = x10 ^ x2 ;
  assign n276 = x26 ^ x18 ;
  assign n301 = n275 & n276 ;
  assign n306 = n302 ^ n301 ;
  assign n273 = x9 ^ x1 ;
  assign n274 = x25 ^ x17 ;
  assign n295 = n273 & n274 ;
  assign n271 = x8 ^ x0 ;
  assign n272 = x24 ^ x16 ;
  assign n294 = n271 & n272 ;
  assign n299 = n295 ^ n294 ;
  assign n320 = n306 ^ n299 ;
  assign n401 = n352 ^ n320 ;
  assign n421 = n413 ^ n401 ;
  assign n422 = n421 ^ n264 ;
  assign n335 = n285 ^ n283 ;
  assign n336 = n286 ^ n284 ;
  assign n337 = n335 & n336 ;
  assign n339 = n337 ^ n333 ;
  assign n328 = n281 ^ n279 ;
  assign n329 = n282 ^ n280 ;
  assign n330 = n328 & n329 ;
  assign n332 = n330 ^ n326 ;
  assign n353 = n339 ^ n332 ;
  assign n303 = n277 ^ n275 ;
  assign n304 = n278 ^ n276 ;
  assign n305 = n303 & n304 ;
  assign n307 = n305 ^ n301 ;
  assign n296 = n273 ^ n271 ;
  assign n297 = n274 ^ n272 ;
  assign n298 = n296 & n297 ;
  assign n300 = n298 ^ n294 ;
  assign n321 = n307 ^ n300 ;
  assign n402 = n353 ^ n321 ;
  assign n423 = n414 ^ n402 ;
  assign n424 = n423 ^ n266 ;
  assign n342 = n285 ^ n281 ;
  assign n343 = n286 ^ n282 ;
  assign n346 = n342 & n343 ;
  assign n340 = n283 ^ n279 ;
  assign n341 = n284 ^ n280 ;
  assign n345 = n340 & n341 ;
  assign n350 = n346 ^ n345 ;
  assign n354 = n352 ^ n350 ;
  assign n355 = n354 ^ n339 ;
  assign n310 = n277 ^ n273 ;
  assign n311 = n278 ^ n274 ;
  assign n314 = n310 & n311 ;
  assign n308 = n275 ^ n271 ;
  assign n309 = n276 ^ n272 ;
  assign n313 = n308 & n309 ;
  assign n318 = n314 ^ n313 ;
  assign n322 = n320 ^ n318 ;
  assign n323 = n322 ^ n307 ;
  assign n403 = n355 ^ n323 ;
  assign n425 = n415 ^ n403 ;
  assign n426 = n425 ^ n268 ;
  assign n347 = n342 ^ n340 ;
  assign n348 = n343 ^ n341 ;
  assign n349 = n347 & n348 ;
  assign n351 = n349 ^ n345 ;
  assign n356 = n353 ^ n351 ;
  assign n344 = n339 ^ n338 ;
  assign n357 = n356 ^ n344 ;
  assign n315 = n310 ^ n308 ;
  assign n316 = n311 ^ n309 ;
  assign n317 = n315 & n316 ;
  assign n319 = n317 ^ n313 ;
  assign n324 = n321 ^ n319 ;
  assign n312 = n307 ^ n306 ;
  assign n325 = n324 ^ n312 ;
  assign n404 = n357 ^ n325 ;
  assign n427 = n416 ^ n404 ;
  assign n428 = n427 ^ n270 ;
  assign n364 = n285 ^ n277 ;
  assign n365 = n286 ^ n278 ;
  assign n377 = n364 & n365 ;
  assign n362 = n283 ^ n275 ;
  assign n363 = n284 ^ n276 ;
  assign n376 = n362 & n363 ;
  assign n381 = n377 ^ n376 ;
  assign n360 = n281 ^ n273 ;
  assign n361 = n282 ^ n274 ;
  assign n370 = n360 & n361 ;
  assign n358 = n279 ^ n271 ;
  assign n359 = n280 ^ n272 ;
  assign n369 = n358 & n359 ;
  assign n374 = n370 ^ n369 ;
  assign n395 = n381 ^ n374 ;
  assign n405 = n401 ^ n395 ;
  assign n406 = n405 ^ n355 ;
  assign n429 = n417 ^ n406 ;
  assign n290 = n268 ^ n259 ;
  assign n430 = n429 ^ n290 ;
  assign n378 = n364 ^ n362 ;
  assign n379 = n365 ^ n363 ;
  assign n380 = n378 & n379 ;
  assign n382 = n380 ^ n376 ;
  assign n371 = n360 ^ n358 ;
  assign n372 = n361 ^ n359 ;
  assign n373 = n371 & n372 ;
  assign n375 = n373 ^ n369 ;
  assign n396 = n382 ^ n375 ;
  assign n407 = n402 ^ n396 ;
  assign n408 = n407 ^ n357 ;
  assign n431 = n418 ^ n408 ;
  assign n291 = n270 ^ n260 ;
  assign n432 = n431 ^ n291 ;
  assign n385 = n364 ^ n360 ;
  assign n386 = n365 ^ n361 ;
  assign n389 = n385 & n386 ;
  assign n383 = n362 ^ n358 ;
  assign n384 = n363 ^ n359 ;
  assign n388 = n383 & n384 ;
  assign n393 = n389 ^ n388 ;
  assign n397 = n395 ^ n393 ;
  assign n398 = n397 ^ n382 ;
  assign n409 = n403 ^ n398 ;
  assign n367 = n357 ^ n352 ;
  assign n410 = n409 ^ n367 ;
  assign n433 = n419 ^ n410 ;
  assign n288 = n270 ^ n264 ;
  assign n292 = n288 ^ n261 ;
  assign n434 = n433 ^ n292 ;
  assign n390 = n385 ^ n383 ;
  assign n391 = n386 ^ n384 ;
  assign n392 = n390 & n391 ;
  assign n394 = n392 ^ n388 ;
  assign n399 = n396 ^ n394 ;
  assign n387 = n382 ^ n381 ;
  assign n400 = n399 ^ n387 ;
  assign n411 = n404 ^ n400 ;
  assign n366 = n357 ^ n355 ;
  assign n368 = n366 ^ n353 ;
  assign n412 = n411 ^ n368 ;
  assign n435 = n420 ^ n412 ;
  assign n287 = n270 ^ n268 ;
  assign n289 = n287 ^ n266 ;
  assign n293 = n289 ^ n262 ;
  assign n436 = n435 ^ n293 ;
  assign y0 = n413 ;
  assign y1 = n414 ;
  assign y2 = n415 ;
  assign y3 = n416 ;
  assign y4 = n417 ;
  assign y5 = n418 ;
  assign y6 = n419 ;
  assign y7 = n420 ;
  assign y8 = n422 ;
  assign y9 = n424 ;
  assign y10 = n426 ;
  assign y11 = n428 ;
  assign y12 = n430 ;
  assign y13 = n432 ;
  assign y14 = n434 ;
  assign y15 = n436 ;
endmodule
