module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 ;
  assign n2120 = x63 & x127 ;
  assign n2119 = x62 & x126 ;
  assign n2124 = n2120 ^ n2119 ;
  assign n2112 = x61 & x125 ;
  assign n2111 = x60 & x124 ;
  assign n2116 = n2112 ^ n2111 ;
  assign n2140 = n2124 ^ n2116 ;
  assign n2085 = x59 & x123 ;
  assign n2084 = x58 & x122 ;
  assign n2089 = n2085 ^ n2084 ;
  assign n2077 = x57 & x121 ;
  assign n2076 = x56 & x120 ;
  assign n2081 = n2077 ^ n2076 ;
  assign n2105 = n2089 ^ n2081 ;
  assign n2192 = n2140 ^ n2105 ;
  assign n1992 = x55 & x119 ;
  assign n1991 = x54 & x118 ;
  assign n1996 = n1992 ^ n1991 ;
  assign n1984 = x53 & x117 ;
  assign n1983 = x52 & x116 ;
  assign n1988 = n1984 ^ n1983 ;
  assign n2012 = n1996 ^ n1988 ;
  assign n1957 = x51 & x115 ;
  assign n1956 = x50 & x114 ;
  assign n1961 = n1957 ^ n1956 ;
  assign n1949 = x49 & x113 ;
  assign n1948 = x48 & x112 ;
  assign n1953 = n1949 ^ n1948 ;
  assign n1977 = n1961 ^ n1953 ;
  assign n2064 = n2012 ^ n1977 ;
  assign n2355 = n2192 ^ n2064 ;
  assign n1689 = x47 & x111 ;
  assign n1688 = x46 & x110 ;
  assign n1693 = n1689 ^ n1688 ;
  assign n1681 = x45 & x109 ;
  assign n1680 = x44 & x108 ;
  assign n1685 = n1681 ^ n1680 ;
  assign n1709 = n1693 ^ n1685 ;
  assign n1654 = x43 & x107 ;
  assign n1653 = x42 & x106 ;
  assign n1658 = n1654 ^ n1653 ;
  assign n1646 = x41 & x105 ;
  assign n1645 = x40 & x104 ;
  assign n1650 = n1646 ^ n1645 ;
  assign n1674 = n1658 ^ n1650 ;
  assign n1761 = n1709 ^ n1674 ;
  assign n1561 = x39 & x103 ;
  assign n1560 = x38 & x102 ;
  assign n1565 = n1561 ^ n1560 ;
  assign n1553 = x37 & x101 ;
  assign n1552 = x36 & x100 ;
  assign n1557 = n1553 ^ n1552 ;
  assign n1581 = n1565 ^ n1557 ;
  assign n1526 = x35 & x99 ;
  assign n1525 = x34 & x98 ;
  assign n1530 = n1526 ^ n1525 ;
  assign n1518 = x33 & x97 ;
  assign n1517 = x32 & x96 ;
  assign n1522 = n1518 ^ n1517 ;
  assign n1546 = n1530 ^ n1522 ;
  assign n1633 = n1581 ^ n1546 ;
  assign n1924 = n1761 ^ n1633 ;
  assign n2857 = n2355 ^ n1924 ;
  assign n732 = x31 & x95 ;
  assign n731 = x30 & x94 ;
  assign n736 = n732 ^ n731 ;
  assign n724 = x29 & x93 ;
  assign n723 = x28 & x92 ;
  assign n728 = n724 ^ n723 ;
  assign n752 = n736 ^ n728 ;
  assign n697 = x27 & x91 ;
  assign n696 = x26 & x90 ;
  assign n701 = n697 ^ n696 ;
  assign n689 = x25 & x89 ;
  assign n688 = x24 & x88 ;
  assign n693 = n689 ^ n688 ;
  assign n717 = n701 ^ n693 ;
  assign n804 = n752 ^ n717 ;
  assign n604 = x23 & x87 ;
  assign n603 = x22 & x86 ;
  assign n608 = n604 ^ n603 ;
  assign n596 = x21 & x85 ;
  assign n595 = x20 & x84 ;
  assign n600 = n596 ^ n595 ;
  assign n624 = n608 ^ n600 ;
  assign n569 = x19 & x83 ;
  assign n568 = x18 & x82 ;
  assign n573 = n569 ^ n568 ;
  assign n561 = x17 & x81 ;
  assign n560 = x16 & x80 ;
  assign n565 = n561 ^ n560 ;
  assign n589 = n573 ^ n565 ;
  assign n676 = n624 ^ n589 ;
  assign n967 = n804 ^ n676 ;
  assign n301 = x15 & x79 ;
  assign n300 = x14 & x78 ;
  assign n305 = n301 ^ n300 ;
  assign n293 = x13 & x77 ;
  assign n292 = x12 & x76 ;
  assign n297 = n293 ^ n292 ;
  assign n321 = n305 ^ n297 ;
  assign n266 = x11 & x75 ;
  assign n265 = x10 & x74 ;
  assign n270 = n266 ^ n265 ;
  assign n258 = x9 & x73 ;
  assign n257 = x8 & x72 ;
  assign n262 = n258 ^ n257 ;
  assign n286 = n270 ^ n262 ;
  assign n373 = n321 ^ n286 ;
  assign n173 = x7 & x71 ;
  assign n172 = x6 & x70 ;
  assign n177 = n173 ^ n172 ;
  assign n165 = x5 & x69 ;
  assign n164 = x4 & x68 ;
  assign n169 = n165 ^ n164 ;
  assign n193 = n177 ^ n169 ;
  assign n138 = x3 & x67 ;
  assign n137 = x2 & x66 ;
  assign n142 = n138 ^ n137 ;
  assign n130 = x1 & x65 ;
  assign n129 = x0 & x64 ;
  assign n134 = n130 ^ n129 ;
  assign n158 = n142 ^ n134 ;
  assign n245 = n193 ^ n158 ;
  assign n536 = n373 ^ n245 ;
  assign n1469 = n967 ^ n536 ;
  assign n4388 = n2857 ^ n1469 ;
  assign n2121 = x63 ^ x62 ;
  assign n2122 = x127 ^ x126 ;
  assign n2123 = n2121 & n2122 ;
  assign n2125 = n2124 ^ n2123 ;
  assign n2126 = n2125 ^ n2120 ;
  assign n2113 = x61 ^ x60 ;
  assign n2114 = x125 ^ x124 ;
  assign n2115 = n2113 & n2114 ;
  assign n2117 = n2116 ^ n2115 ;
  assign n2118 = n2117 ^ n2112 ;
  assign n2141 = n2126 ^ n2118 ;
  assign n2086 = x59 ^ x58 ;
  assign n2087 = x123 ^ x122 ;
  assign n2088 = n2086 & n2087 ;
  assign n2090 = n2089 ^ n2088 ;
  assign n2091 = n2090 ^ n2085 ;
  assign n2078 = x57 ^ x56 ;
  assign n2079 = x121 ^ x120 ;
  assign n2080 = n2078 & n2079 ;
  assign n2082 = n2081 ^ n2080 ;
  assign n2083 = n2082 ^ n2077 ;
  assign n2106 = n2091 ^ n2083 ;
  assign n2193 = n2141 ^ n2106 ;
  assign n1993 = x55 ^ x54 ;
  assign n1994 = x119 ^ x118 ;
  assign n1995 = n1993 & n1994 ;
  assign n1997 = n1996 ^ n1995 ;
  assign n1998 = n1997 ^ n1992 ;
  assign n1985 = x53 ^ x52 ;
  assign n1986 = x117 ^ x116 ;
  assign n1987 = n1985 & n1986 ;
  assign n1989 = n1988 ^ n1987 ;
  assign n1990 = n1989 ^ n1984 ;
  assign n2013 = n1998 ^ n1990 ;
  assign n1958 = x51 ^ x50 ;
  assign n1959 = x115 ^ x114 ;
  assign n1960 = n1958 & n1959 ;
  assign n1962 = n1961 ^ n1960 ;
  assign n1963 = n1962 ^ n1957 ;
  assign n1950 = x49 ^ x48 ;
  assign n1951 = x113 ^ x112 ;
  assign n1952 = n1950 & n1951 ;
  assign n1954 = n1953 ^ n1952 ;
  assign n1955 = n1954 ^ n1949 ;
  assign n1978 = n1963 ^ n1955 ;
  assign n2065 = n2013 ^ n1978 ;
  assign n2356 = n2193 ^ n2065 ;
  assign n1690 = x47 ^ x46 ;
  assign n1691 = x111 ^ x110 ;
  assign n1692 = n1690 & n1691 ;
  assign n1694 = n1693 ^ n1692 ;
  assign n1695 = n1694 ^ n1689 ;
  assign n1682 = x45 ^ x44 ;
  assign n1683 = x109 ^ x108 ;
  assign n1684 = n1682 & n1683 ;
  assign n1686 = n1685 ^ n1684 ;
  assign n1687 = n1686 ^ n1681 ;
  assign n1710 = n1695 ^ n1687 ;
  assign n1655 = x43 ^ x42 ;
  assign n1656 = x107 ^ x106 ;
  assign n1657 = n1655 & n1656 ;
  assign n1659 = n1658 ^ n1657 ;
  assign n1660 = n1659 ^ n1654 ;
  assign n1647 = x41 ^ x40 ;
  assign n1648 = x105 ^ x104 ;
  assign n1649 = n1647 & n1648 ;
  assign n1651 = n1650 ^ n1649 ;
  assign n1652 = n1651 ^ n1646 ;
  assign n1675 = n1660 ^ n1652 ;
  assign n1762 = n1710 ^ n1675 ;
  assign n1562 = x39 ^ x38 ;
  assign n1563 = x103 ^ x102 ;
  assign n1564 = n1562 & n1563 ;
  assign n1566 = n1565 ^ n1564 ;
  assign n1567 = n1566 ^ n1561 ;
  assign n1554 = x37 ^ x36 ;
  assign n1555 = x101 ^ x100 ;
  assign n1556 = n1554 & n1555 ;
  assign n1558 = n1557 ^ n1556 ;
  assign n1559 = n1558 ^ n1553 ;
  assign n1582 = n1567 ^ n1559 ;
  assign n1527 = x35 ^ x34 ;
  assign n1528 = x99 ^ x98 ;
  assign n1529 = n1527 & n1528 ;
  assign n1531 = n1530 ^ n1529 ;
  assign n1532 = n1531 ^ n1526 ;
  assign n1519 = x33 ^ x32 ;
  assign n1520 = x97 ^ x96 ;
  assign n1521 = n1519 & n1520 ;
  assign n1523 = n1522 ^ n1521 ;
  assign n1524 = n1523 ^ n1518 ;
  assign n1547 = n1532 ^ n1524 ;
  assign n1634 = n1582 ^ n1547 ;
  assign n1925 = n1762 ^ n1634 ;
  assign n2858 = n2356 ^ n1925 ;
  assign n733 = x31 ^ x30 ;
  assign n734 = x95 ^ x94 ;
  assign n735 = n733 & n734 ;
  assign n737 = n736 ^ n735 ;
  assign n738 = n737 ^ n732 ;
  assign n725 = x29 ^ x28 ;
  assign n726 = x93 ^ x92 ;
  assign n727 = n725 & n726 ;
  assign n729 = n728 ^ n727 ;
  assign n730 = n729 ^ n724 ;
  assign n753 = n738 ^ n730 ;
  assign n698 = x27 ^ x26 ;
  assign n699 = x91 ^ x90 ;
  assign n700 = n698 & n699 ;
  assign n702 = n701 ^ n700 ;
  assign n703 = n702 ^ n697 ;
  assign n690 = x25 ^ x24 ;
  assign n691 = x89 ^ x88 ;
  assign n692 = n690 & n691 ;
  assign n694 = n693 ^ n692 ;
  assign n695 = n694 ^ n689 ;
  assign n718 = n703 ^ n695 ;
  assign n805 = n753 ^ n718 ;
  assign n605 = x23 ^ x22 ;
  assign n606 = x87 ^ x86 ;
  assign n607 = n605 & n606 ;
  assign n609 = n608 ^ n607 ;
  assign n610 = n609 ^ n604 ;
  assign n597 = x21 ^ x20 ;
  assign n598 = x85 ^ x84 ;
  assign n599 = n597 & n598 ;
  assign n601 = n600 ^ n599 ;
  assign n602 = n601 ^ n596 ;
  assign n625 = n610 ^ n602 ;
  assign n570 = x19 ^ x18 ;
  assign n571 = x83 ^ x82 ;
  assign n572 = n570 & n571 ;
  assign n574 = n573 ^ n572 ;
  assign n575 = n574 ^ n569 ;
  assign n562 = x17 ^ x16 ;
  assign n563 = x81 ^ x80 ;
  assign n564 = n562 & n563 ;
  assign n566 = n565 ^ n564 ;
  assign n567 = n566 ^ n561 ;
  assign n590 = n575 ^ n567 ;
  assign n677 = n625 ^ n590 ;
  assign n968 = n805 ^ n677 ;
  assign n302 = x15 ^ x14 ;
  assign n303 = x79 ^ x78 ;
  assign n304 = n302 & n303 ;
  assign n306 = n305 ^ n304 ;
  assign n307 = n306 ^ n301 ;
  assign n294 = x13 ^ x12 ;
  assign n295 = x77 ^ x76 ;
  assign n296 = n294 & n295 ;
  assign n298 = n297 ^ n296 ;
  assign n299 = n298 ^ n293 ;
  assign n322 = n307 ^ n299 ;
  assign n267 = x11 ^ x10 ;
  assign n268 = x75 ^ x74 ;
  assign n269 = n267 & n268 ;
  assign n271 = n270 ^ n269 ;
  assign n272 = n271 ^ n266 ;
  assign n259 = x9 ^ x8 ;
  assign n260 = x73 ^ x72 ;
  assign n261 = n259 & n260 ;
  assign n263 = n262 ^ n261 ;
  assign n264 = n263 ^ n258 ;
  assign n287 = n272 ^ n264 ;
  assign n374 = n322 ^ n287 ;
  assign n174 = x7 ^ x6 ;
  assign n175 = x71 ^ x70 ;
  assign n176 = n174 & n175 ;
  assign n178 = n177 ^ n176 ;
  assign n179 = n178 ^ n173 ;
  assign n166 = x5 ^ x4 ;
  assign n167 = x69 ^ x68 ;
  assign n168 = n166 & n167 ;
  assign n170 = n169 ^ n168 ;
  assign n171 = n170 ^ n165 ;
  assign n194 = n179 ^ n171 ;
  assign n139 = x3 ^ x2 ;
  assign n140 = x67 ^ x66 ;
  assign n141 = n139 & n140 ;
  assign n143 = n142 ^ n141 ;
  assign n144 = n143 ^ n138 ;
  assign n131 = x1 ^ x0 ;
  assign n132 = x65 ^ x64 ;
  assign n133 = n131 & n132 ;
  assign n135 = n134 ^ n133 ;
  assign n136 = n135 ^ n130 ;
  assign n159 = n144 ^ n136 ;
  assign n246 = n194 ^ n159 ;
  assign n537 = n374 ^ n246 ;
  assign n1470 = n968 ^ n537 ;
  assign n4389 = n2858 ^ n1470 ;
  assign n2130 = x63 ^ x61 ;
  assign n2131 = x127 ^ x125 ;
  assign n2133 = n2130 & n2131 ;
  assign n2128 = x62 ^ x60 ;
  assign n2129 = x126 ^ x124 ;
  assign n2132 = n2128 & n2129 ;
  assign n2137 = n2133 ^ n2132 ;
  assign n2142 = n2140 ^ n2137 ;
  assign n2143 = n2142 ^ n2126 ;
  assign n2095 = x59 ^ x57 ;
  assign n2096 = x123 ^ x121 ;
  assign n2098 = n2095 & n2096 ;
  assign n2093 = x58 ^ x56 ;
  assign n2094 = x122 ^ x120 ;
  assign n2097 = n2093 & n2094 ;
  assign n2102 = n2098 ^ n2097 ;
  assign n2107 = n2105 ^ n2102 ;
  assign n2108 = n2107 ^ n2091 ;
  assign n2194 = n2143 ^ n2108 ;
  assign n2002 = x55 ^ x53 ;
  assign n2003 = x119 ^ x117 ;
  assign n2005 = n2002 & n2003 ;
  assign n2000 = x54 ^ x52 ;
  assign n2001 = x118 ^ x116 ;
  assign n2004 = n2000 & n2001 ;
  assign n2009 = n2005 ^ n2004 ;
  assign n2014 = n2012 ^ n2009 ;
  assign n2015 = n2014 ^ n1998 ;
  assign n1967 = x51 ^ x49 ;
  assign n1968 = x115 ^ x113 ;
  assign n1970 = n1967 & n1968 ;
  assign n1965 = x50 ^ x48 ;
  assign n1966 = x114 ^ x112 ;
  assign n1969 = n1965 & n1966 ;
  assign n1974 = n1970 ^ n1969 ;
  assign n1979 = n1977 ^ n1974 ;
  assign n1980 = n1979 ^ n1963 ;
  assign n2066 = n2015 ^ n1980 ;
  assign n2357 = n2194 ^ n2066 ;
  assign n1699 = x47 ^ x45 ;
  assign n1700 = x111 ^ x109 ;
  assign n1702 = n1699 & n1700 ;
  assign n1697 = x46 ^ x44 ;
  assign n1698 = x110 ^ x108 ;
  assign n1701 = n1697 & n1698 ;
  assign n1706 = n1702 ^ n1701 ;
  assign n1711 = n1709 ^ n1706 ;
  assign n1712 = n1711 ^ n1695 ;
  assign n1664 = x43 ^ x41 ;
  assign n1665 = x107 ^ x105 ;
  assign n1667 = n1664 & n1665 ;
  assign n1662 = x42 ^ x40 ;
  assign n1663 = x106 ^ x104 ;
  assign n1666 = n1662 & n1663 ;
  assign n1671 = n1667 ^ n1666 ;
  assign n1676 = n1674 ^ n1671 ;
  assign n1677 = n1676 ^ n1660 ;
  assign n1763 = n1712 ^ n1677 ;
  assign n1571 = x39 ^ x37 ;
  assign n1572 = x103 ^ x101 ;
  assign n1574 = n1571 & n1572 ;
  assign n1569 = x38 ^ x36 ;
  assign n1570 = x102 ^ x100 ;
  assign n1573 = n1569 & n1570 ;
  assign n1578 = n1574 ^ n1573 ;
  assign n1583 = n1581 ^ n1578 ;
  assign n1584 = n1583 ^ n1567 ;
  assign n1536 = x35 ^ x33 ;
  assign n1537 = x99 ^ x97 ;
  assign n1539 = n1536 & n1537 ;
  assign n1534 = x34 ^ x32 ;
  assign n1535 = x98 ^ x96 ;
  assign n1538 = n1534 & n1535 ;
  assign n1543 = n1539 ^ n1538 ;
  assign n1548 = n1546 ^ n1543 ;
  assign n1549 = n1548 ^ n1532 ;
  assign n1635 = n1584 ^ n1549 ;
  assign n1926 = n1763 ^ n1635 ;
  assign n2859 = n2357 ^ n1926 ;
  assign n742 = x31 ^ x29 ;
  assign n743 = x95 ^ x93 ;
  assign n745 = n742 & n743 ;
  assign n740 = x30 ^ x28 ;
  assign n741 = x94 ^ x92 ;
  assign n744 = n740 & n741 ;
  assign n749 = n745 ^ n744 ;
  assign n754 = n752 ^ n749 ;
  assign n755 = n754 ^ n738 ;
  assign n707 = x27 ^ x25 ;
  assign n708 = x91 ^ x89 ;
  assign n710 = n707 & n708 ;
  assign n705 = x26 ^ x24 ;
  assign n706 = x90 ^ x88 ;
  assign n709 = n705 & n706 ;
  assign n714 = n710 ^ n709 ;
  assign n719 = n717 ^ n714 ;
  assign n720 = n719 ^ n703 ;
  assign n806 = n755 ^ n720 ;
  assign n614 = x23 ^ x21 ;
  assign n615 = x87 ^ x85 ;
  assign n617 = n614 & n615 ;
  assign n612 = x22 ^ x20 ;
  assign n613 = x86 ^ x84 ;
  assign n616 = n612 & n613 ;
  assign n621 = n617 ^ n616 ;
  assign n626 = n624 ^ n621 ;
  assign n627 = n626 ^ n610 ;
  assign n579 = x19 ^ x17 ;
  assign n580 = x83 ^ x81 ;
  assign n582 = n579 & n580 ;
  assign n577 = x18 ^ x16 ;
  assign n578 = x82 ^ x80 ;
  assign n581 = n577 & n578 ;
  assign n586 = n582 ^ n581 ;
  assign n591 = n589 ^ n586 ;
  assign n592 = n591 ^ n575 ;
  assign n678 = n627 ^ n592 ;
  assign n969 = n806 ^ n678 ;
  assign n311 = x15 ^ x13 ;
  assign n312 = x79 ^ x77 ;
  assign n314 = n311 & n312 ;
  assign n309 = x14 ^ x12 ;
  assign n310 = x78 ^ x76 ;
  assign n313 = n309 & n310 ;
  assign n318 = n314 ^ n313 ;
  assign n323 = n321 ^ n318 ;
  assign n324 = n323 ^ n307 ;
  assign n276 = x11 ^ x9 ;
  assign n277 = x75 ^ x73 ;
  assign n279 = n276 & n277 ;
  assign n274 = x10 ^ x8 ;
  assign n275 = x74 ^ x72 ;
  assign n278 = n274 & n275 ;
  assign n283 = n279 ^ n278 ;
  assign n288 = n286 ^ n283 ;
  assign n289 = n288 ^ n272 ;
  assign n375 = n324 ^ n289 ;
  assign n183 = x7 ^ x5 ;
  assign n184 = x71 ^ x69 ;
  assign n186 = n183 & n184 ;
  assign n181 = x6 ^ x4 ;
  assign n182 = x70 ^ x68 ;
  assign n185 = n181 & n182 ;
  assign n190 = n186 ^ n185 ;
  assign n195 = n193 ^ n190 ;
  assign n196 = n195 ^ n179 ;
  assign n148 = x3 ^ x1 ;
  assign n149 = x67 ^ x65 ;
  assign n151 = n148 & n149 ;
  assign n146 = x2 ^ x0 ;
  assign n147 = x66 ^ x64 ;
  assign n150 = n146 & n147 ;
  assign n155 = n151 ^ n150 ;
  assign n160 = n158 ^ n155 ;
  assign n161 = n160 ^ n144 ;
  assign n247 = n196 ^ n161 ;
  assign n538 = n375 ^ n247 ;
  assign n1471 = n969 ^ n538 ;
  assign n4390 = n2859 ^ n1471 ;
  assign n2134 = n2130 ^ n2128 ;
  assign n2135 = n2131 ^ n2129 ;
  assign n2136 = n2134 & n2135 ;
  assign n2138 = n2137 ^ n2136 ;
  assign n2139 = n2138 ^ n2133 ;
  assign n2144 = n2141 ^ n2139 ;
  assign n2127 = n2126 ^ n2124 ;
  assign n2145 = n2144 ^ n2127 ;
  assign n2099 = n2095 ^ n2093 ;
  assign n2100 = n2096 ^ n2094 ;
  assign n2101 = n2099 & n2100 ;
  assign n2103 = n2102 ^ n2101 ;
  assign n2104 = n2103 ^ n2098 ;
  assign n2109 = n2106 ^ n2104 ;
  assign n2092 = n2091 ^ n2089 ;
  assign n2110 = n2109 ^ n2092 ;
  assign n2195 = n2145 ^ n2110 ;
  assign n2006 = n2002 ^ n2000 ;
  assign n2007 = n2003 ^ n2001 ;
  assign n2008 = n2006 & n2007 ;
  assign n2010 = n2009 ^ n2008 ;
  assign n2011 = n2010 ^ n2005 ;
  assign n2016 = n2013 ^ n2011 ;
  assign n1999 = n1998 ^ n1996 ;
  assign n2017 = n2016 ^ n1999 ;
  assign n1971 = n1967 ^ n1965 ;
  assign n1972 = n1968 ^ n1966 ;
  assign n1973 = n1971 & n1972 ;
  assign n1975 = n1974 ^ n1973 ;
  assign n1976 = n1975 ^ n1970 ;
  assign n1981 = n1978 ^ n1976 ;
  assign n1964 = n1963 ^ n1961 ;
  assign n1982 = n1981 ^ n1964 ;
  assign n2067 = n2017 ^ n1982 ;
  assign n2358 = n2195 ^ n2067 ;
  assign n1703 = n1699 ^ n1697 ;
  assign n1704 = n1700 ^ n1698 ;
  assign n1705 = n1703 & n1704 ;
  assign n1707 = n1706 ^ n1705 ;
  assign n1708 = n1707 ^ n1702 ;
  assign n1713 = n1710 ^ n1708 ;
  assign n1696 = n1695 ^ n1693 ;
  assign n1714 = n1713 ^ n1696 ;
  assign n1668 = n1664 ^ n1662 ;
  assign n1669 = n1665 ^ n1663 ;
  assign n1670 = n1668 & n1669 ;
  assign n1672 = n1671 ^ n1670 ;
  assign n1673 = n1672 ^ n1667 ;
  assign n1678 = n1675 ^ n1673 ;
  assign n1661 = n1660 ^ n1658 ;
  assign n1679 = n1678 ^ n1661 ;
  assign n1764 = n1714 ^ n1679 ;
  assign n1575 = n1571 ^ n1569 ;
  assign n1576 = n1572 ^ n1570 ;
  assign n1577 = n1575 & n1576 ;
  assign n1579 = n1578 ^ n1577 ;
  assign n1580 = n1579 ^ n1574 ;
  assign n1585 = n1582 ^ n1580 ;
  assign n1568 = n1567 ^ n1565 ;
  assign n1586 = n1585 ^ n1568 ;
  assign n1540 = n1536 ^ n1534 ;
  assign n1541 = n1537 ^ n1535 ;
  assign n1542 = n1540 & n1541 ;
  assign n1544 = n1543 ^ n1542 ;
  assign n1545 = n1544 ^ n1539 ;
  assign n1550 = n1547 ^ n1545 ;
  assign n1533 = n1532 ^ n1530 ;
  assign n1551 = n1550 ^ n1533 ;
  assign n1636 = n1586 ^ n1551 ;
  assign n1927 = n1764 ^ n1636 ;
  assign n2860 = n2358 ^ n1927 ;
  assign n746 = n742 ^ n740 ;
  assign n747 = n743 ^ n741 ;
  assign n748 = n746 & n747 ;
  assign n750 = n749 ^ n748 ;
  assign n751 = n750 ^ n745 ;
  assign n756 = n753 ^ n751 ;
  assign n739 = n738 ^ n736 ;
  assign n757 = n756 ^ n739 ;
  assign n711 = n707 ^ n705 ;
  assign n712 = n708 ^ n706 ;
  assign n713 = n711 & n712 ;
  assign n715 = n714 ^ n713 ;
  assign n716 = n715 ^ n710 ;
  assign n721 = n718 ^ n716 ;
  assign n704 = n703 ^ n701 ;
  assign n722 = n721 ^ n704 ;
  assign n807 = n757 ^ n722 ;
  assign n618 = n614 ^ n612 ;
  assign n619 = n615 ^ n613 ;
  assign n620 = n618 & n619 ;
  assign n622 = n621 ^ n620 ;
  assign n623 = n622 ^ n617 ;
  assign n628 = n625 ^ n623 ;
  assign n611 = n610 ^ n608 ;
  assign n629 = n628 ^ n611 ;
  assign n583 = n579 ^ n577 ;
  assign n584 = n580 ^ n578 ;
  assign n585 = n583 & n584 ;
  assign n587 = n586 ^ n585 ;
  assign n588 = n587 ^ n582 ;
  assign n593 = n590 ^ n588 ;
  assign n576 = n575 ^ n573 ;
  assign n594 = n593 ^ n576 ;
  assign n679 = n629 ^ n594 ;
  assign n970 = n807 ^ n679 ;
  assign n315 = n311 ^ n309 ;
  assign n316 = n312 ^ n310 ;
  assign n317 = n315 & n316 ;
  assign n319 = n318 ^ n317 ;
  assign n320 = n319 ^ n314 ;
  assign n325 = n322 ^ n320 ;
  assign n308 = n307 ^ n305 ;
  assign n326 = n325 ^ n308 ;
  assign n280 = n276 ^ n274 ;
  assign n281 = n277 ^ n275 ;
  assign n282 = n280 & n281 ;
  assign n284 = n283 ^ n282 ;
  assign n285 = n284 ^ n279 ;
  assign n290 = n287 ^ n285 ;
  assign n273 = n272 ^ n270 ;
  assign n291 = n290 ^ n273 ;
  assign n376 = n326 ^ n291 ;
  assign n187 = n183 ^ n181 ;
  assign n188 = n184 ^ n182 ;
  assign n189 = n187 & n188 ;
  assign n191 = n190 ^ n189 ;
  assign n192 = n191 ^ n186 ;
  assign n197 = n194 ^ n192 ;
  assign n180 = n179 ^ n177 ;
  assign n198 = n197 ^ n180 ;
  assign n152 = n148 ^ n146 ;
  assign n153 = n149 ^ n147 ;
  assign n154 = n152 & n153 ;
  assign n156 = n155 ^ n154 ;
  assign n157 = n156 ^ n151 ;
  assign n162 = n159 ^ n157 ;
  assign n145 = n144 ^ n142 ;
  assign n163 = n162 ^ n145 ;
  assign n248 = n198 ^ n163 ;
  assign n539 = n376 ^ n248 ;
  assign n1472 = n970 ^ n539 ;
  assign n4391 = n2860 ^ n1472 ;
  assign n2155 = x63 ^ x59 ;
  assign n2156 = x127 ^ x123 ;
  assign n2166 = n2155 & n2156 ;
  assign n2153 = x62 ^ x58 ;
  assign n2154 = x126 ^ x122 ;
  assign n2165 = n2153 & n2154 ;
  assign n2170 = n2166 ^ n2165 ;
  assign n2151 = x61 ^ x57 ;
  assign n2152 = x125 ^ x121 ;
  assign n2158 = n2151 & n2152 ;
  assign n2149 = x60 ^ x56 ;
  assign n2150 = x124 ^ x120 ;
  assign n2157 = n2149 & n2150 ;
  assign n2162 = n2158 ^ n2157 ;
  assign n2186 = n2170 ^ n2162 ;
  assign n2196 = n2192 ^ n2186 ;
  assign n2197 = n2196 ^ n2143 ;
  assign n2027 = x55 ^ x51 ;
  assign n2028 = x119 ^ x115 ;
  assign n2038 = n2027 & n2028 ;
  assign n2025 = x54 ^ x50 ;
  assign n2026 = x118 ^ x114 ;
  assign n2037 = n2025 & n2026 ;
  assign n2042 = n2038 ^ n2037 ;
  assign n2023 = x53 ^ x49 ;
  assign n2024 = x117 ^ x113 ;
  assign n2030 = n2023 & n2024 ;
  assign n2021 = x52 ^ x48 ;
  assign n2022 = x116 ^ x112 ;
  assign n2029 = n2021 & n2022 ;
  assign n2034 = n2030 ^ n2029 ;
  assign n2058 = n2042 ^ n2034 ;
  assign n2068 = n2064 ^ n2058 ;
  assign n2069 = n2068 ^ n2015 ;
  assign n2359 = n2197 ^ n2069 ;
  assign n1724 = x47 ^ x43 ;
  assign n1725 = x111 ^ x107 ;
  assign n1735 = n1724 & n1725 ;
  assign n1722 = x46 ^ x42 ;
  assign n1723 = x110 ^ x106 ;
  assign n1734 = n1722 & n1723 ;
  assign n1739 = n1735 ^ n1734 ;
  assign n1720 = x45 ^ x41 ;
  assign n1721 = x109 ^ x105 ;
  assign n1727 = n1720 & n1721 ;
  assign n1718 = x44 ^ x40 ;
  assign n1719 = x108 ^ x104 ;
  assign n1726 = n1718 & n1719 ;
  assign n1731 = n1727 ^ n1726 ;
  assign n1755 = n1739 ^ n1731 ;
  assign n1765 = n1761 ^ n1755 ;
  assign n1766 = n1765 ^ n1712 ;
  assign n1596 = x39 ^ x35 ;
  assign n1597 = x103 ^ x99 ;
  assign n1607 = n1596 & n1597 ;
  assign n1594 = x38 ^ x34 ;
  assign n1595 = x102 ^ x98 ;
  assign n1606 = n1594 & n1595 ;
  assign n1611 = n1607 ^ n1606 ;
  assign n1592 = x37 ^ x33 ;
  assign n1593 = x101 ^ x97 ;
  assign n1599 = n1592 & n1593 ;
  assign n1590 = x36 ^ x32 ;
  assign n1591 = x100 ^ x96 ;
  assign n1598 = n1590 & n1591 ;
  assign n1603 = n1599 ^ n1598 ;
  assign n1627 = n1611 ^ n1603 ;
  assign n1637 = n1633 ^ n1627 ;
  assign n1638 = n1637 ^ n1584 ;
  assign n1928 = n1766 ^ n1638 ;
  assign n2861 = n2359 ^ n1928 ;
  assign n767 = x31 ^ x27 ;
  assign n768 = x95 ^ x91 ;
  assign n778 = n767 & n768 ;
  assign n765 = x30 ^ x26 ;
  assign n766 = x94 ^ x90 ;
  assign n777 = n765 & n766 ;
  assign n782 = n778 ^ n777 ;
  assign n763 = x29 ^ x25 ;
  assign n764 = x93 ^ x89 ;
  assign n770 = n763 & n764 ;
  assign n761 = x28 ^ x24 ;
  assign n762 = x92 ^ x88 ;
  assign n769 = n761 & n762 ;
  assign n774 = n770 ^ n769 ;
  assign n798 = n782 ^ n774 ;
  assign n808 = n804 ^ n798 ;
  assign n809 = n808 ^ n755 ;
  assign n639 = x23 ^ x19 ;
  assign n640 = x87 ^ x83 ;
  assign n650 = n639 & n640 ;
  assign n637 = x22 ^ x18 ;
  assign n638 = x86 ^ x82 ;
  assign n649 = n637 & n638 ;
  assign n654 = n650 ^ n649 ;
  assign n635 = x21 ^ x17 ;
  assign n636 = x85 ^ x81 ;
  assign n642 = n635 & n636 ;
  assign n633 = x20 ^ x16 ;
  assign n634 = x84 ^ x80 ;
  assign n641 = n633 & n634 ;
  assign n646 = n642 ^ n641 ;
  assign n670 = n654 ^ n646 ;
  assign n680 = n676 ^ n670 ;
  assign n681 = n680 ^ n627 ;
  assign n971 = n809 ^ n681 ;
  assign n336 = x15 ^ x11 ;
  assign n337 = x79 ^ x75 ;
  assign n347 = n336 & n337 ;
  assign n334 = x14 ^ x10 ;
  assign n335 = x78 ^ x74 ;
  assign n346 = n334 & n335 ;
  assign n351 = n347 ^ n346 ;
  assign n332 = x13 ^ x9 ;
  assign n333 = x77 ^ x73 ;
  assign n339 = n332 & n333 ;
  assign n330 = x12 ^ x8 ;
  assign n331 = x76 ^ x72 ;
  assign n338 = n330 & n331 ;
  assign n343 = n339 ^ n338 ;
  assign n367 = n351 ^ n343 ;
  assign n377 = n373 ^ n367 ;
  assign n378 = n377 ^ n324 ;
  assign n208 = x7 ^ x3 ;
  assign n209 = x71 ^ x67 ;
  assign n219 = n208 & n209 ;
  assign n206 = x6 ^ x2 ;
  assign n207 = x70 ^ x66 ;
  assign n218 = n206 & n207 ;
  assign n223 = n219 ^ n218 ;
  assign n204 = x5 ^ x1 ;
  assign n205 = x69 ^ x65 ;
  assign n211 = n204 & n205 ;
  assign n202 = x4 ^ x0 ;
  assign n203 = x68 ^ x64 ;
  assign n210 = n202 & n203 ;
  assign n215 = n211 ^ n210 ;
  assign n239 = n223 ^ n215 ;
  assign n249 = n245 ^ n239 ;
  assign n250 = n249 ^ n196 ;
  assign n540 = n378 ^ n250 ;
  assign n1473 = n971 ^ n540 ;
  assign n4392 = n2861 ^ n1473 ;
  assign n2167 = n2155 ^ n2153 ;
  assign n2168 = n2156 ^ n2154 ;
  assign n2169 = n2167 & n2168 ;
  assign n2171 = n2170 ^ n2169 ;
  assign n2172 = n2171 ^ n2166 ;
  assign n2159 = n2151 ^ n2149 ;
  assign n2160 = n2152 ^ n2150 ;
  assign n2161 = n2159 & n2160 ;
  assign n2163 = n2162 ^ n2161 ;
  assign n2164 = n2163 ^ n2158 ;
  assign n2187 = n2172 ^ n2164 ;
  assign n2198 = n2193 ^ n2187 ;
  assign n2199 = n2198 ^ n2145 ;
  assign n2039 = n2027 ^ n2025 ;
  assign n2040 = n2028 ^ n2026 ;
  assign n2041 = n2039 & n2040 ;
  assign n2043 = n2042 ^ n2041 ;
  assign n2044 = n2043 ^ n2038 ;
  assign n2031 = n2023 ^ n2021 ;
  assign n2032 = n2024 ^ n2022 ;
  assign n2033 = n2031 & n2032 ;
  assign n2035 = n2034 ^ n2033 ;
  assign n2036 = n2035 ^ n2030 ;
  assign n2059 = n2044 ^ n2036 ;
  assign n2070 = n2065 ^ n2059 ;
  assign n2071 = n2070 ^ n2017 ;
  assign n2360 = n2199 ^ n2071 ;
  assign n1736 = n1724 ^ n1722 ;
  assign n1737 = n1725 ^ n1723 ;
  assign n1738 = n1736 & n1737 ;
  assign n1740 = n1739 ^ n1738 ;
  assign n1741 = n1740 ^ n1735 ;
  assign n1728 = n1720 ^ n1718 ;
  assign n1729 = n1721 ^ n1719 ;
  assign n1730 = n1728 & n1729 ;
  assign n1732 = n1731 ^ n1730 ;
  assign n1733 = n1732 ^ n1727 ;
  assign n1756 = n1741 ^ n1733 ;
  assign n1767 = n1762 ^ n1756 ;
  assign n1768 = n1767 ^ n1714 ;
  assign n1608 = n1596 ^ n1594 ;
  assign n1609 = n1597 ^ n1595 ;
  assign n1610 = n1608 & n1609 ;
  assign n1612 = n1611 ^ n1610 ;
  assign n1613 = n1612 ^ n1607 ;
  assign n1600 = n1592 ^ n1590 ;
  assign n1601 = n1593 ^ n1591 ;
  assign n1602 = n1600 & n1601 ;
  assign n1604 = n1603 ^ n1602 ;
  assign n1605 = n1604 ^ n1599 ;
  assign n1628 = n1613 ^ n1605 ;
  assign n1639 = n1634 ^ n1628 ;
  assign n1640 = n1639 ^ n1586 ;
  assign n1929 = n1768 ^ n1640 ;
  assign n2862 = n2360 ^ n1929 ;
  assign n779 = n767 ^ n765 ;
  assign n780 = n768 ^ n766 ;
  assign n781 = n779 & n780 ;
  assign n783 = n782 ^ n781 ;
  assign n784 = n783 ^ n778 ;
  assign n771 = n763 ^ n761 ;
  assign n772 = n764 ^ n762 ;
  assign n773 = n771 & n772 ;
  assign n775 = n774 ^ n773 ;
  assign n776 = n775 ^ n770 ;
  assign n799 = n784 ^ n776 ;
  assign n810 = n805 ^ n799 ;
  assign n811 = n810 ^ n757 ;
  assign n651 = n639 ^ n637 ;
  assign n652 = n640 ^ n638 ;
  assign n653 = n651 & n652 ;
  assign n655 = n654 ^ n653 ;
  assign n656 = n655 ^ n650 ;
  assign n643 = n635 ^ n633 ;
  assign n644 = n636 ^ n634 ;
  assign n645 = n643 & n644 ;
  assign n647 = n646 ^ n645 ;
  assign n648 = n647 ^ n642 ;
  assign n671 = n656 ^ n648 ;
  assign n682 = n677 ^ n671 ;
  assign n683 = n682 ^ n629 ;
  assign n972 = n811 ^ n683 ;
  assign n348 = n336 ^ n334 ;
  assign n349 = n337 ^ n335 ;
  assign n350 = n348 & n349 ;
  assign n352 = n351 ^ n350 ;
  assign n353 = n352 ^ n347 ;
  assign n340 = n332 ^ n330 ;
  assign n341 = n333 ^ n331 ;
  assign n342 = n340 & n341 ;
  assign n344 = n343 ^ n342 ;
  assign n345 = n344 ^ n339 ;
  assign n368 = n353 ^ n345 ;
  assign n379 = n374 ^ n368 ;
  assign n380 = n379 ^ n326 ;
  assign n220 = n208 ^ n206 ;
  assign n221 = n209 ^ n207 ;
  assign n222 = n220 & n221 ;
  assign n224 = n223 ^ n222 ;
  assign n225 = n224 ^ n219 ;
  assign n212 = n204 ^ n202 ;
  assign n213 = n205 ^ n203 ;
  assign n214 = n212 & n213 ;
  assign n216 = n215 ^ n214 ;
  assign n217 = n216 ^ n211 ;
  assign n240 = n225 ^ n217 ;
  assign n251 = n246 ^ n240 ;
  assign n252 = n251 ^ n198 ;
  assign n541 = n380 ^ n252 ;
  assign n1474 = n972 ^ n541 ;
  assign n4393 = n2862 ^ n1474 ;
  assign n2176 = n2155 ^ n2151 ;
  assign n2177 = n2156 ^ n2152 ;
  assign n2179 = n2176 & n2177 ;
  assign n2174 = n2153 ^ n2149 ;
  assign n2175 = n2154 ^ n2150 ;
  assign n2178 = n2174 & n2175 ;
  assign n2183 = n2179 ^ n2178 ;
  assign n2188 = n2186 ^ n2183 ;
  assign n2189 = n2188 ^ n2172 ;
  assign n2200 = n2194 ^ n2189 ;
  assign n2147 = n2145 ^ n2140 ;
  assign n2201 = n2200 ^ n2147 ;
  assign n2048 = n2027 ^ n2023 ;
  assign n2049 = n2028 ^ n2024 ;
  assign n2051 = n2048 & n2049 ;
  assign n2046 = n2025 ^ n2021 ;
  assign n2047 = n2026 ^ n2022 ;
  assign n2050 = n2046 & n2047 ;
  assign n2055 = n2051 ^ n2050 ;
  assign n2060 = n2058 ^ n2055 ;
  assign n2061 = n2060 ^ n2044 ;
  assign n2072 = n2066 ^ n2061 ;
  assign n2019 = n2017 ^ n2012 ;
  assign n2073 = n2072 ^ n2019 ;
  assign n2361 = n2201 ^ n2073 ;
  assign n1745 = n1724 ^ n1720 ;
  assign n1746 = n1725 ^ n1721 ;
  assign n1748 = n1745 & n1746 ;
  assign n1743 = n1722 ^ n1718 ;
  assign n1744 = n1723 ^ n1719 ;
  assign n1747 = n1743 & n1744 ;
  assign n1752 = n1748 ^ n1747 ;
  assign n1757 = n1755 ^ n1752 ;
  assign n1758 = n1757 ^ n1741 ;
  assign n1769 = n1763 ^ n1758 ;
  assign n1716 = n1714 ^ n1709 ;
  assign n1770 = n1769 ^ n1716 ;
  assign n1617 = n1596 ^ n1592 ;
  assign n1618 = n1597 ^ n1593 ;
  assign n1620 = n1617 & n1618 ;
  assign n1615 = n1594 ^ n1590 ;
  assign n1616 = n1595 ^ n1591 ;
  assign n1619 = n1615 & n1616 ;
  assign n1624 = n1620 ^ n1619 ;
  assign n1629 = n1627 ^ n1624 ;
  assign n1630 = n1629 ^ n1613 ;
  assign n1641 = n1635 ^ n1630 ;
  assign n1588 = n1586 ^ n1581 ;
  assign n1642 = n1641 ^ n1588 ;
  assign n1930 = n1770 ^ n1642 ;
  assign n2863 = n2361 ^ n1930 ;
  assign n788 = n767 ^ n763 ;
  assign n789 = n768 ^ n764 ;
  assign n791 = n788 & n789 ;
  assign n786 = n765 ^ n761 ;
  assign n787 = n766 ^ n762 ;
  assign n790 = n786 & n787 ;
  assign n795 = n791 ^ n790 ;
  assign n800 = n798 ^ n795 ;
  assign n801 = n800 ^ n784 ;
  assign n812 = n806 ^ n801 ;
  assign n759 = n757 ^ n752 ;
  assign n813 = n812 ^ n759 ;
  assign n660 = n639 ^ n635 ;
  assign n661 = n640 ^ n636 ;
  assign n663 = n660 & n661 ;
  assign n658 = n637 ^ n633 ;
  assign n659 = n638 ^ n634 ;
  assign n662 = n658 & n659 ;
  assign n667 = n663 ^ n662 ;
  assign n672 = n670 ^ n667 ;
  assign n673 = n672 ^ n656 ;
  assign n684 = n678 ^ n673 ;
  assign n631 = n629 ^ n624 ;
  assign n685 = n684 ^ n631 ;
  assign n973 = n813 ^ n685 ;
  assign n357 = n336 ^ n332 ;
  assign n358 = n337 ^ n333 ;
  assign n360 = n357 & n358 ;
  assign n355 = n334 ^ n330 ;
  assign n356 = n335 ^ n331 ;
  assign n359 = n355 & n356 ;
  assign n364 = n360 ^ n359 ;
  assign n369 = n367 ^ n364 ;
  assign n370 = n369 ^ n353 ;
  assign n381 = n375 ^ n370 ;
  assign n328 = n326 ^ n321 ;
  assign n382 = n381 ^ n328 ;
  assign n229 = n208 ^ n204 ;
  assign n230 = n209 ^ n205 ;
  assign n232 = n229 & n230 ;
  assign n227 = n206 ^ n202 ;
  assign n228 = n207 ^ n203 ;
  assign n231 = n227 & n228 ;
  assign n236 = n232 ^ n231 ;
  assign n241 = n239 ^ n236 ;
  assign n242 = n241 ^ n225 ;
  assign n253 = n247 ^ n242 ;
  assign n200 = n198 ^ n193 ;
  assign n254 = n253 ^ n200 ;
  assign n542 = n382 ^ n254 ;
  assign n1475 = n973 ^ n542 ;
  assign n4394 = n2863 ^ n1475 ;
  assign n2180 = n2176 ^ n2174 ;
  assign n2181 = n2177 ^ n2175 ;
  assign n2182 = n2180 & n2181 ;
  assign n2184 = n2183 ^ n2182 ;
  assign n2185 = n2184 ^ n2179 ;
  assign n2190 = n2187 ^ n2185 ;
  assign n2173 = n2172 ^ n2170 ;
  assign n2191 = n2190 ^ n2173 ;
  assign n2202 = n2195 ^ n2191 ;
  assign n2146 = n2145 ^ n2143 ;
  assign n2148 = n2146 ^ n2141 ;
  assign n2203 = n2202 ^ n2148 ;
  assign n2052 = n2048 ^ n2046 ;
  assign n2053 = n2049 ^ n2047 ;
  assign n2054 = n2052 & n2053 ;
  assign n2056 = n2055 ^ n2054 ;
  assign n2057 = n2056 ^ n2051 ;
  assign n2062 = n2059 ^ n2057 ;
  assign n2045 = n2044 ^ n2042 ;
  assign n2063 = n2062 ^ n2045 ;
  assign n2074 = n2067 ^ n2063 ;
  assign n2018 = n2017 ^ n2015 ;
  assign n2020 = n2018 ^ n2013 ;
  assign n2075 = n2074 ^ n2020 ;
  assign n2362 = n2203 ^ n2075 ;
  assign n1749 = n1745 ^ n1743 ;
  assign n1750 = n1746 ^ n1744 ;
  assign n1751 = n1749 & n1750 ;
  assign n1753 = n1752 ^ n1751 ;
  assign n1754 = n1753 ^ n1748 ;
  assign n1759 = n1756 ^ n1754 ;
  assign n1742 = n1741 ^ n1739 ;
  assign n1760 = n1759 ^ n1742 ;
  assign n1771 = n1764 ^ n1760 ;
  assign n1715 = n1714 ^ n1712 ;
  assign n1717 = n1715 ^ n1710 ;
  assign n1772 = n1771 ^ n1717 ;
  assign n1621 = n1617 ^ n1615 ;
  assign n1622 = n1618 ^ n1616 ;
  assign n1623 = n1621 & n1622 ;
  assign n1625 = n1624 ^ n1623 ;
  assign n1626 = n1625 ^ n1620 ;
  assign n1631 = n1628 ^ n1626 ;
  assign n1614 = n1613 ^ n1611 ;
  assign n1632 = n1631 ^ n1614 ;
  assign n1643 = n1636 ^ n1632 ;
  assign n1587 = n1586 ^ n1584 ;
  assign n1589 = n1587 ^ n1582 ;
  assign n1644 = n1643 ^ n1589 ;
  assign n1931 = n1772 ^ n1644 ;
  assign n2864 = n2362 ^ n1931 ;
  assign n792 = n788 ^ n786 ;
  assign n793 = n789 ^ n787 ;
  assign n794 = n792 & n793 ;
  assign n796 = n795 ^ n794 ;
  assign n797 = n796 ^ n791 ;
  assign n802 = n799 ^ n797 ;
  assign n785 = n784 ^ n782 ;
  assign n803 = n802 ^ n785 ;
  assign n814 = n807 ^ n803 ;
  assign n758 = n757 ^ n755 ;
  assign n760 = n758 ^ n753 ;
  assign n815 = n814 ^ n760 ;
  assign n664 = n660 ^ n658 ;
  assign n665 = n661 ^ n659 ;
  assign n666 = n664 & n665 ;
  assign n668 = n667 ^ n666 ;
  assign n669 = n668 ^ n663 ;
  assign n674 = n671 ^ n669 ;
  assign n657 = n656 ^ n654 ;
  assign n675 = n674 ^ n657 ;
  assign n686 = n679 ^ n675 ;
  assign n630 = n629 ^ n627 ;
  assign n632 = n630 ^ n625 ;
  assign n687 = n686 ^ n632 ;
  assign n974 = n815 ^ n687 ;
  assign n361 = n357 ^ n355 ;
  assign n362 = n358 ^ n356 ;
  assign n363 = n361 & n362 ;
  assign n365 = n364 ^ n363 ;
  assign n366 = n365 ^ n360 ;
  assign n371 = n368 ^ n366 ;
  assign n354 = n353 ^ n351 ;
  assign n372 = n371 ^ n354 ;
  assign n383 = n376 ^ n372 ;
  assign n327 = n326 ^ n324 ;
  assign n329 = n327 ^ n322 ;
  assign n384 = n383 ^ n329 ;
  assign n233 = n229 ^ n227 ;
  assign n234 = n230 ^ n228 ;
  assign n235 = n233 & n234 ;
  assign n237 = n236 ^ n235 ;
  assign n238 = n237 ^ n232 ;
  assign n243 = n240 ^ n238 ;
  assign n226 = n225 ^ n223 ;
  assign n244 = n243 ^ n226 ;
  assign n255 = n248 ^ n244 ;
  assign n199 = n198 ^ n196 ;
  assign n201 = n199 ^ n194 ;
  assign n256 = n255 ^ n201 ;
  assign n543 = n384 ^ n256 ;
  assign n1476 = n974 ^ n543 ;
  assign n4395 = n2864 ^ n1476 ;
  assign n2225 = x63 ^ x55 ;
  assign n2226 = x127 ^ x119 ;
  assign n2271 = n2225 & n2226 ;
  assign n2223 = x62 ^ x54 ;
  assign n2224 = x126 ^ x118 ;
  assign n2270 = n2223 & n2224 ;
  assign n2275 = n2271 ^ n2270 ;
  assign n2221 = x61 ^ x53 ;
  assign n2222 = x125 ^ x117 ;
  assign n2263 = n2221 & n2222 ;
  assign n2219 = x60 ^ x52 ;
  assign n2220 = x124 ^ x116 ;
  assign n2262 = n2219 & n2220 ;
  assign n2267 = n2263 ^ n2262 ;
  assign n2291 = n2275 ^ n2267 ;
  assign n2217 = x59 ^ x51 ;
  assign n2218 = x123 ^ x115 ;
  assign n2236 = n2217 & n2218 ;
  assign n2215 = x58 ^ x50 ;
  assign n2216 = x122 ^ x114 ;
  assign n2235 = n2215 & n2216 ;
  assign n2240 = n2236 ^ n2235 ;
  assign n2213 = x57 ^ x49 ;
  assign n2214 = x121 ^ x113 ;
  assign n2228 = n2213 & n2214 ;
  assign n2211 = x56 ^ x48 ;
  assign n2212 = x120 ^ x112 ;
  assign n2227 = n2211 & n2212 ;
  assign n2232 = n2228 ^ n2227 ;
  assign n2256 = n2240 ^ n2232 ;
  assign n2343 = n2291 ^ n2256 ;
  assign n2363 = n2355 ^ n2343 ;
  assign n2364 = n2363 ^ n2197 ;
  assign n1794 = x47 ^ x39 ;
  assign n1795 = x111 ^ x103 ;
  assign n1840 = n1794 & n1795 ;
  assign n1792 = x46 ^ x38 ;
  assign n1793 = x110 ^ x102 ;
  assign n1839 = n1792 & n1793 ;
  assign n1844 = n1840 ^ n1839 ;
  assign n1790 = x45 ^ x37 ;
  assign n1791 = x109 ^ x101 ;
  assign n1832 = n1790 & n1791 ;
  assign n1788 = x44 ^ x36 ;
  assign n1789 = x108 ^ x100 ;
  assign n1831 = n1788 & n1789 ;
  assign n1836 = n1832 ^ n1831 ;
  assign n1860 = n1844 ^ n1836 ;
  assign n1786 = x43 ^ x35 ;
  assign n1787 = x107 ^ x99 ;
  assign n1805 = n1786 & n1787 ;
  assign n1784 = x42 ^ x34 ;
  assign n1785 = x106 ^ x98 ;
  assign n1804 = n1784 & n1785 ;
  assign n1809 = n1805 ^ n1804 ;
  assign n1782 = x41 ^ x33 ;
  assign n1783 = x105 ^ x97 ;
  assign n1797 = n1782 & n1783 ;
  assign n1780 = x40 ^ x32 ;
  assign n1781 = x104 ^ x96 ;
  assign n1796 = n1780 & n1781 ;
  assign n1801 = n1797 ^ n1796 ;
  assign n1825 = n1809 ^ n1801 ;
  assign n1912 = n1860 ^ n1825 ;
  assign n1932 = n1924 ^ n1912 ;
  assign n1933 = n1932 ^ n1766 ;
  assign n2865 = n2364 ^ n1933 ;
  assign n837 = x31 ^ x23 ;
  assign n838 = x95 ^ x87 ;
  assign n883 = n837 & n838 ;
  assign n835 = x30 ^ x22 ;
  assign n836 = x94 ^ x86 ;
  assign n882 = n835 & n836 ;
  assign n887 = n883 ^ n882 ;
  assign n833 = x29 ^ x21 ;
  assign n834 = x93 ^ x85 ;
  assign n875 = n833 & n834 ;
  assign n831 = x28 ^ x20 ;
  assign n832 = x92 ^ x84 ;
  assign n874 = n831 & n832 ;
  assign n879 = n875 ^ n874 ;
  assign n903 = n887 ^ n879 ;
  assign n829 = x27 ^ x19 ;
  assign n830 = x91 ^ x83 ;
  assign n848 = n829 & n830 ;
  assign n827 = x26 ^ x18 ;
  assign n828 = x90 ^ x82 ;
  assign n847 = n827 & n828 ;
  assign n852 = n848 ^ n847 ;
  assign n825 = x25 ^ x17 ;
  assign n826 = x89 ^ x81 ;
  assign n840 = n825 & n826 ;
  assign n823 = x24 ^ x16 ;
  assign n824 = x88 ^ x80 ;
  assign n839 = n823 & n824 ;
  assign n844 = n840 ^ n839 ;
  assign n868 = n852 ^ n844 ;
  assign n955 = n903 ^ n868 ;
  assign n975 = n967 ^ n955 ;
  assign n976 = n975 ^ n809 ;
  assign n406 = x15 ^ x7 ;
  assign n407 = x79 ^ x71 ;
  assign n452 = n406 & n407 ;
  assign n404 = x14 ^ x6 ;
  assign n405 = x78 ^ x70 ;
  assign n451 = n404 & n405 ;
  assign n456 = n452 ^ n451 ;
  assign n402 = x13 ^ x5 ;
  assign n403 = x77 ^ x69 ;
  assign n444 = n402 & n403 ;
  assign n400 = x12 ^ x4 ;
  assign n401 = x76 ^ x68 ;
  assign n443 = n400 & n401 ;
  assign n448 = n444 ^ n443 ;
  assign n472 = n456 ^ n448 ;
  assign n398 = x11 ^ x3 ;
  assign n399 = x75 ^ x67 ;
  assign n417 = n398 & n399 ;
  assign n396 = x10 ^ x2 ;
  assign n397 = x74 ^ x66 ;
  assign n416 = n396 & n397 ;
  assign n421 = n417 ^ n416 ;
  assign n394 = x9 ^ x1 ;
  assign n395 = x73 ^ x65 ;
  assign n409 = n394 & n395 ;
  assign n392 = x8 ^ x0 ;
  assign n393 = x72 ^ x64 ;
  assign n408 = n392 & n393 ;
  assign n413 = n409 ^ n408 ;
  assign n437 = n421 ^ n413 ;
  assign n524 = n472 ^ n437 ;
  assign n544 = n536 ^ n524 ;
  assign n545 = n544 ^ n378 ;
  assign n1477 = n976 ^ n545 ;
  assign n4396 = n2865 ^ n1477 ;
  assign n2272 = n2225 ^ n2223 ;
  assign n2273 = n2226 ^ n2224 ;
  assign n2274 = n2272 & n2273 ;
  assign n2276 = n2275 ^ n2274 ;
  assign n2277 = n2276 ^ n2271 ;
  assign n2264 = n2221 ^ n2219 ;
  assign n2265 = n2222 ^ n2220 ;
  assign n2266 = n2264 & n2265 ;
  assign n2268 = n2267 ^ n2266 ;
  assign n2269 = n2268 ^ n2263 ;
  assign n2292 = n2277 ^ n2269 ;
  assign n2237 = n2217 ^ n2215 ;
  assign n2238 = n2218 ^ n2216 ;
  assign n2239 = n2237 & n2238 ;
  assign n2241 = n2240 ^ n2239 ;
  assign n2242 = n2241 ^ n2236 ;
  assign n2229 = n2213 ^ n2211 ;
  assign n2230 = n2214 ^ n2212 ;
  assign n2231 = n2229 & n2230 ;
  assign n2233 = n2232 ^ n2231 ;
  assign n2234 = n2233 ^ n2228 ;
  assign n2257 = n2242 ^ n2234 ;
  assign n2344 = n2292 ^ n2257 ;
  assign n2365 = n2356 ^ n2344 ;
  assign n2366 = n2365 ^ n2199 ;
  assign n1841 = n1794 ^ n1792 ;
  assign n1842 = n1795 ^ n1793 ;
  assign n1843 = n1841 & n1842 ;
  assign n1845 = n1844 ^ n1843 ;
  assign n1846 = n1845 ^ n1840 ;
  assign n1833 = n1790 ^ n1788 ;
  assign n1834 = n1791 ^ n1789 ;
  assign n1835 = n1833 & n1834 ;
  assign n1837 = n1836 ^ n1835 ;
  assign n1838 = n1837 ^ n1832 ;
  assign n1861 = n1846 ^ n1838 ;
  assign n1806 = n1786 ^ n1784 ;
  assign n1807 = n1787 ^ n1785 ;
  assign n1808 = n1806 & n1807 ;
  assign n1810 = n1809 ^ n1808 ;
  assign n1811 = n1810 ^ n1805 ;
  assign n1798 = n1782 ^ n1780 ;
  assign n1799 = n1783 ^ n1781 ;
  assign n1800 = n1798 & n1799 ;
  assign n1802 = n1801 ^ n1800 ;
  assign n1803 = n1802 ^ n1797 ;
  assign n1826 = n1811 ^ n1803 ;
  assign n1913 = n1861 ^ n1826 ;
  assign n1934 = n1925 ^ n1913 ;
  assign n1935 = n1934 ^ n1768 ;
  assign n2866 = n2366 ^ n1935 ;
  assign n884 = n837 ^ n835 ;
  assign n885 = n838 ^ n836 ;
  assign n886 = n884 & n885 ;
  assign n888 = n887 ^ n886 ;
  assign n889 = n888 ^ n883 ;
  assign n876 = n833 ^ n831 ;
  assign n877 = n834 ^ n832 ;
  assign n878 = n876 & n877 ;
  assign n880 = n879 ^ n878 ;
  assign n881 = n880 ^ n875 ;
  assign n904 = n889 ^ n881 ;
  assign n849 = n829 ^ n827 ;
  assign n850 = n830 ^ n828 ;
  assign n851 = n849 & n850 ;
  assign n853 = n852 ^ n851 ;
  assign n854 = n853 ^ n848 ;
  assign n841 = n825 ^ n823 ;
  assign n842 = n826 ^ n824 ;
  assign n843 = n841 & n842 ;
  assign n845 = n844 ^ n843 ;
  assign n846 = n845 ^ n840 ;
  assign n869 = n854 ^ n846 ;
  assign n956 = n904 ^ n869 ;
  assign n977 = n968 ^ n956 ;
  assign n978 = n977 ^ n811 ;
  assign n453 = n406 ^ n404 ;
  assign n454 = n407 ^ n405 ;
  assign n455 = n453 & n454 ;
  assign n457 = n456 ^ n455 ;
  assign n458 = n457 ^ n452 ;
  assign n445 = n402 ^ n400 ;
  assign n446 = n403 ^ n401 ;
  assign n447 = n445 & n446 ;
  assign n449 = n448 ^ n447 ;
  assign n450 = n449 ^ n444 ;
  assign n473 = n458 ^ n450 ;
  assign n418 = n398 ^ n396 ;
  assign n419 = n399 ^ n397 ;
  assign n420 = n418 & n419 ;
  assign n422 = n421 ^ n420 ;
  assign n423 = n422 ^ n417 ;
  assign n410 = n394 ^ n392 ;
  assign n411 = n395 ^ n393 ;
  assign n412 = n410 & n411 ;
  assign n414 = n413 ^ n412 ;
  assign n415 = n414 ^ n409 ;
  assign n438 = n423 ^ n415 ;
  assign n525 = n473 ^ n438 ;
  assign n546 = n537 ^ n525 ;
  assign n547 = n546 ^ n380 ;
  assign n1478 = n978 ^ n547 ;
  assign n4397 = n2866 ^ n1478 ;
  assign n2281 = n2225 ^ n2221 ;
  assign n2282 = n2226 ^ n2222 ;
  assign n2284 = n2281 & n2282 ;
  assign n2279 = n2223 ^ n2219 ;
  assign n2280 = n2224 ^ n2220 ;
  assign n2283 = n2279 & n2280 ;
  assign n2288 = n2284 ^ n2283 ;
  assign n2293 = n2291 ^ n2288 ;
  assign n2294 = n2293 ^ n2277 ;
  assign n2246 = n2217 ^ n2213 ;
  assign n2247 = n2218 ^ n2214 ;
  assign n2249 = n2246 & n2247 ;
  assign n2244 = n2215 ^ n2211 ;
  assign n2245 = n2216 ^ n2212 ;
  assign n2248 = n2244 & n2245 ;
  assign n2253 = n2249 ^ n2248 ;
  assign n2258 = n2256 ^ n2253 ;
  assign n2259 = n2258 ^ n2242 ;
  assign n2345 = n2294 ^ n2259 ;
  assign n2367 = n2357 ^ n2345 ;
  assign n2368 = n2367 ^ n2201 ;
  assign n1850 = n1794 ^ n1790 ;
  assign n1851 = n1795 ^ n1791 ;
  assign n1853 = n1850 & n1851 ;
  assign n1848 = n1792 ^ n1788 ;
  assign n1849 = n1793 ^ n1789 ;
  assign n1852 = n1848 & n1849 ;
  assign n1857 = n1853 ^ n1852 ;
  assign n1862 = n1860 ^ n1857 ;
  assign n1863 = n1862 ^ n1846 ;
  assign n1815 = n1786 ^ n1782 ;
  assign n1816 = n1787 ^ n1783 ;
  assign n1818 = n1815 & n1816 ;
  assign n1813 = n1784 ^ n1780 ;
  assign n1814 = n1785 ^ n1781 ;
  assign n1817 = n1813 & n1814 ;
  assign n1822 = n1818 ^ n1817 ;
  assign n1827 = n1825 ^ n1822 ;
  assign n1828 = n1827 ^ n1811 ;
  assign n1914 = n1863 ^ n1828 ;
  assign n1936 = n1926 ^ n1914 ;
  assign n1937 = n1936 ^ n1770 ;
  assign n2867 = n2368 ^ n1937 ;
  assign n893 = n837 ^ n833 ;
  assign n894 = n838 ^ n834 ;
  assign n896 = n893 & n894 ;
  assign n891 = n835 ^ n831 ;
  assign n892 = n836 ^ n832 ;
  assign n895 = n891 & n892 ;
  assign n900 = n896 ^ n895 ;
  assign n905 = n903 ^ n900 ;
  assign n906 = n905 ^ n889 ;
  assign n858 = n829 ^ n825 ;
  assign n859 = n830 ^ n826 ;
  assign n861 = n858 & n859 ;
  assign n856 = n827 ^ n823 ;
  assign n857 = n828 ^ n824 ;
  assign n860 = n856 & n857 ;
  assign n865 = n861 ^ n860 ;
  assign n870 = n868 ^ n865 ;
  assign n871 = n870 ^ n854 ;
  assign n957 = n906 ^ n871 ;
  assign n979 = n969 ^ n957 ;
  assign n980 = n979 ^ n813 ;
  assign n462 = n406 ^ n402 ;
  assign n463 = n407 ^ n403 ;
  assign n465 = n462 & n463 ;
  assign n460 = n404 ^ n400 ;
  assign n461 = n405 ^ n401 ;
  assign n464 = n460 & n461 ;
  assign n469 = n465 ^ n464 ;
  assign n474 = n472 ^ n469 ;
  assign n475 = n474 ^ n458 ;
  assign n427 = n398 ^ n394 ;
  assign n428 = n399 ^ n395 ;
  assign n430 = n427 & n428 ;
  assign n425 = n396 ^ n392 ;
  assign n426 = n397 ^ n393 ;
  assign n429 = n425 & n426 ;
  assign n434 = n430 ^ n429 ;
  assign n439 = n437 ^ n434 ;
  assign n440 = n439 ^ n423 ;
  assign n526 = n475 ^ n440 ;
  assign n548 = n538 ^ n526 ;
  assign n549 = n548 ^ n382 ;
  assign n1479 = n980 ^ n549 ;
  assign n4398 = n2867 ^ n1479 ;
  assign n2285 = n2281 ^ n2279 ;
  assign n2286 = n2282 ^ n2280 ;
  assign n2287 = n2285 & n2286 ;
  assign n2289 = n2288 ^ n2287 ;
  assign n2290 = n2289 ^ n2284 ;
  assign n2295 = n2292 ^ n2290 ;
  assign n2278 = n2277 ^ n2275 ;
  assign n2296 = n2295 ^ n2278 ;
  assign n2250 = n2246 ^ n2244 ;
  assign n2251 = n2247 ^ n2245 ;
  assign n2252 = n2250 & n2251 ;
  assign n2254 = n2253 ^ n2252 ;
  assign n2255 = n2254 ^ n2249 ;
  assign n2260 = n2257 ^ n2255 ;
  assign n2243 = n2242 ^ n2240 ;
  assign n2261 = n2260 ^ n2243 ;
  assign n2346 = n2296 ^ n2261 ;
  assign n2369 = n2358 ^ n2346 ;
  assign n2370 = n2369 ^ n2203 ;
  assign n1854 = n1850 ^ n1848 ;
  assign n1855 = n1851 ^ n1849 ;
  assign n1856 = n1854 & n1855 ;
  assign n1858 = n1857 ^ n1856 ;
  assign n1859 = n1858 ^ n1853 ;
  assign n1864 = n1861 ^ n1859 ;
  assign n1847 = n1846 ^ n1844 ;
  assign n1865 = n1864 ^ n1847 ;
  assign n1819 = n1815 ^ n1813 ;
  assign n1820 = n1816 ^ n1814 ;
  assign n1821 = n1819 & n1820 ;
  assign n1823 = n1822 ^ n1821 ;
  assign n1824 = n1823 ^ n1818 ;
  assign n1829 = n1826 ^ n1824 ;
  assign n1812 = n1811 ^ n1809 ;
  assign n1830 = n1829 ^ n1812 ;
  assign n1915 = n1865 ^ n1830 ;
  assign n1938 = n1927 ^ n1915 ;
  assign n1939 = n1938 ^ n1772 ;
  assign n2868 = n2370 ^ n1939 ;
  assign n897 = n893 ^ n891 ;
  assign n898 = n894 ^ n892 ;
  assign n899 = n897 & n898 ;
  assign n901 = n900 ^ n899 ;
  assign n902 = n901 ^ n896 ;
  assign n907 = n904 ^ n902 ;
  assign n890 = n889 ^ n887 ;
  assign n908 = n907 ^ n890 ;
  assign n862 = n858 ^ n856 ;
  assign n863 = n859 ^ n857 ;
  assign n864 = n862 & n863 ;
  assign n866 = n865 ^ n864 ;
  assign n867 = n866 ^ n861 ;
  assign n872 = n869 ^ n867 ;
  assign n855 = n854 ^ n852 ;
  assign n873 = n872 ^ n855 ;
  assign n958 = n908 ^ n873 ;
  assign n981 = n970 ^ n958 ;
  assign n982 = n981 ^ n815 ;
  assign n466 = n462 ^ n460 ;
  assign n467 = n463 ^ n461 ;
  assign n468 = n466 & n467 ;
  assign n470 = n469 ^ n468 ;
  assign n471 = n470 ^ n465 ;
  assign n476 = n473 ^ n471 ;
  assign n459 = n458 ^ n456 ;
  assign n477 = n476 ^ n459 ;
  assign n431 = n427 ^ n425 ;
  assign n432 = n428 ^ n426 ;
  assign n433 = n431 & n432 ;
  assign n435 = n434 ^ n433 ;
  assign n436 = n435 ^ n430 ;
  assign n441 = n438 ^ n436 ;
  assign n424 = n423 ^ n421 ;
  assign n442 = n441 ^ n424 ;
  assign n527 = n477 ^ n442 ;
  assign n550 = n539 ^ n527 ;
  assign n551 = n550 ^ n384 ;
  assign n1480 = n982 ^ n551 ;
  assign n4399 = n2868 ^ n1480 ;
  assign n2306 = n2225 ^ n2217 ;
  assign n2307 = n2226 ^ n2218 ;
  assign n2317 = n2306 & n2307 ;
  assign n2304 = n2223 ^ n2215 ;
  assign n2305 = n2224 ^ n2216 ;
  assign n2316 = n2304 & n2305 ;
  assign n2321 = n2317 ^ n2316 ;
  assign n2302 = n2221 ^ n2213 ;
  assign n2303 = n2222 ^ n2214 ;
  assign n2309 = n2302 & n2303 ;
  assign n2300 = n2219 ^ n2211 ;
  assign n2301 = n2220 ^ n2212 ;
  assign n2308 = n2300 & n2301 ;
  assign n2313 = n2309 ^ n2308 ;
  assign n2337 = n2321 ^ n2313 ;
  assign n2347 = n2343 ^ n2337 ;
  assign n2348 = n2347 ^ n2294 ;
  assign n2371 = n2359 ^ n2348 ;
  assign n2207 = n2201 ^ n2192 ;
  assign n2372 = n2371 ^ n2207 ;
  assign n1875 = n1794 ^ n1786 ;
  assign n1876 = n1795 ^ n1787 ;
  assign n1886 = n1875 & n1876 ;
  assign n1873 = n1792 ^ n1784 ;
  assign n1874 = n1793 ^ n1785 ;
  assign n1885 = n1873 & n1874 ;
  assign n1890 = n1886 ^ n1885 ;
  assign n1871 = n1790 ^ n1782 ;
  assign n1872 = n1791 ^ n1783 ;
  assign n1878 = n1871 & n1872 ;
  assign n1869 = n1788 ^ n1780 ;
  assign n1870 = n1789 ^ n1781 ;
  assign n1877 = n1869 & n1870 ;
  assign n1882 = n1878 ^ n1877 ;
  assign n1906 = n1890 ^ n1882 ;
  assign n1916 = n1912 ^ n1906 ;
  assign n1917 = n1916 ^ n1863 ;
  assign n1940 = n1928 ^ n1917 ;
  assign n1776 = n1770 ^ n1761 ;
  assign n1941 = n1940 ^ n1776 ;
  assign n2869 = n2372 ^ n1941 ;
  assign n918 = n837 ^ n829 ;
  assign n919 = n838 ^ n830 ;
  assign n929 = n918 & n919 ;
  assign n916 = n835 ^ n827 ;
  assign n917 = n836 ^ n828 ;
  assign n928 = n916 & n917 ;
  assign n933 = n929 ^ n928 ;
  assign n914 = n833 ^ n825 ;
  assign n915 = n834 ^ n826 ;
  assign n921 = n914 & n915 ;
  assign n912 = n831 ^ n823 ;
  assign n913 = n832 ^ n824 ;
  assign n920 = n912 & n913 ;
  assign n925 = n921 ^ n920 ;
  assign n949 = n933 ^ n925 ;
  assign n959 = n955 ^ n949 ;
  assign n960 = n959 ^ n906 ;
  assign n983 = n971 ^ n960 ;
  assign n819 = n813 ^ n804 ;
  assign n984 = n983 ^ n819 ;
  assign n487 = n406 ^ n398 ;
  assign n488 = n407 ^ n399 ;
  assign n498 = n487 & n488 ;
  assign n485 = n404 ^ n396 ;
  assign n486 = n405 ^ n397 ;
  assign n497 = n485 & n486 ;
  assign n502 = n498 ^ n497 ;
  assign n483 = n402 ^ n394 ;
  assign n484 = n403 ^ n395 ;
  assign n490 = n483 & n484 ;
  assign n481 = n400 ^ n392 ;
  assign n482 = n401 ^ n393 ;
  assign n489 = n481 & n482 ;
  assign n494 = n490 ^ n489 ;
  assign n518 = n502 ^ n494 ;
  assign n528 = n524 ^ n518 ;
  assign n529 = n528 ^ n475 ;
  assign n552 = n540 ^ n529 ;
  assign n388 = n382 ^ n373 ;
  assign n553 = n552 ^ n388 ;
  assign n1481 = n984 ^ n553 ;
  assign n4400 = n2869 ^ n1481 ;
  assign n2318 = n2306 ^ n2304 ;
  assign n2319 = n2307 ^ n2305 ;
  assign n2320 = n2318 & n2319 ;
  assign n2322 = n2321 ^ n2320 ;
  assign n2323 = n2322 ^ n2317 ;
  assign n2310 = n2302 ^ n2300 ;
  assign n2311 = n2303 ^ n2301 ;
  assign n2312 = n2310 & n2311 ;
  assign n2314 = n2313 ^ n2312 ;
  assign n2315 = n2314 ^ n2309 ;
  assign n2338 = n2323 ^ n2315 ;
  assign n2349 = n2344 ^ n2338 ;
  assign n2350 = n2349 ^ n2296 ;
  assign n2373 = n2360 ^ n2350 ;
  assign n2208 = n2203 ^ n2193 ;
  assign n2374 = n2373 ^ n2208 ;
  assign n1887 = n1875 ^ n1873 ;
  assign n1888 = n1876 ^ n1874 ;
  assign n1889 = n1887 & n1888 ;
  assign n1891 = n1890 ^ n1889 ;
  assign n1892 = n1891 ^ n1886 ;
  assign n1879 = n1871 ^ n1869 ;
  assign n1880 = n1872 ^ n1870 ;
  assign n1881 = n1879 & n1880 ;
  assign n1883 = n1882 ^ n1881 ;
  assign n1884 = n1883 ^ n1878 ;
  assign n1907 = n1892 ^ n1884 ;
  assign n1918 = n1913 ^ n1907 ;
  assign n1919 = n1918 ^ n1865 ;
  assign n1942 = n1929 ^ n1919 ;
  assign n1777 = n1772 ^ n1762 ;
  assign n1943 = n1942 ^ n1777 ;
  assign n2870 = n2374 ^ n1943 ;
  assign n930 = n918 ^ n916 ;
  assign n931 = n919 ^ n917 ;
  assign n932 = n930 & n931 ;
  assign n934 = n933 ^ n932 ;
  assign n935 = n934 ^ n929 ;
  assign n922 = n914 ^ n912 ;
  assign n923 = n915 ^ n913 ;
  assign n924 = n922 & n923 ;
  assign n926 = n925 ^ n924 ;
  assign n927 = n926 ^ n921 ;
  assign n950 = n935 ^ n927 ;
  assign n961 = n956 ^ n950 ;
  assign n962 = n961 ^ n908 ;
  assign n985 = n972 ^ n962 ;
  assign n820 = n815 ^ n805 ;
  assign n986 = n985 ^ n820 ;
  assign n499 = n487 ^ n485 ;
  assign n500 = n488 ^ n486 ;
  assign n501 = n499 & n500 ;
  assign n503 = n502 ^ n501 ;
  assign n504 = n503 ^ n498 ;
  assign n491 = n483 ^ n481 ;
  assign n492 = n484 ^ n482 ;
  assign n493 = n491 & n492 ;
  assign n495 = n494 ^ n493 ;
  assign n496 = n495 ^ n490 ;
  assign n519 = n504 ^ n496 ;
  assign n530 = n525 ^ n519 ;
  assign n531 = n530 ^ n477 ;
  assign n554 = n541 ^ n531 ;
  assign n389 = n384 ^ n374 ;
  assign n555 = n554 ^ n389 ;
  assign n1482 = n986 ^ n555 ;
  assign n4401 = n2870 ^ n1482 ;
  assign n2327 = n2306 ^ n2302 ;
  assign n2328 = n2307 ^ n2303 ;
  assign n2330 = n2327 & n2328 ;
  assign n2325 = n2304 ^ n2300 ;
  assign n2326 = n2305 ^ n2301 ;
  assign n2329 = n2325 & n2326 ;
  assign n2334 = n2330 ^ n2329 ;
  assign n2339 = n2337 ^ n2334 ;
  assign n2340 = n2339 ^ n2323 ;
  assign n2351 = n2345 ^ n2340 ;
  assign n2298 = n2296 ^ n2291 ;
  assign n2352 = n2351 ^ n2298 ;
  assign n2375 = n2361 ^ n2352 ;
  assign n2205 = n2203 ^ n2197 ;
  assign n2209 = n2205 ^ n2194 ;
  assign n2376 = n2375 ^ n2209 ;
  assign n1896 = n1875 ^ n1871 ;
  assign n1897 = n1876 ^ n1872 ;
  assign n1899 = n1896 & n1897 ;
  assign n1894 = n1873 ^ n1869 ;
  assign n1895 = n1874 ^ n1870 ;
  assign n1898 = n1894 & n1895 ;
  assign n1903 = n1899 ^ n1898 ;
  assign n1908 = n1906 ^ n1903 ;
  assign n1909 = n1908 ^ n1892 ;
  assign n1920 = n1914 ^ n1909 ;
  assign n1867 = n1865 ^ n1860 ;
  assign n1921 = n1920 ^ n1867 ;
  assign n1944 = n1930 ^ n1921 ;
  assign n1774 = n1772 ^ n1766 ;
  assign n1778 = n1774 ^ n1763 ;
  assign n1945 = n1944 ^ n1778 ;
  assign n2871 = n2376 ^ n1945 ;
  assign n939 = n918 ^ n914 ;
  assign n940 = n919 ^ n915 ;
  assign n942 = n939 & n940 ;
  assign n937 = n916 ^ n912 ;
  assign n938 = n917 ^ n913 ;
  assign n941 = n937 & n938 ;
  assign n946 = n942 ^ n941 ;
  assign n951 = n949 ^ n946 ;
  assign n952 = n951 ^ n935 ;
  assign n963 = n957 ^ n952 ;
  assign n910 = n908 ^ n903 ;
  assign n964 = n963 ^ n910 ;
  assign n987 = n973 ^ n964 ;
  assign n817 = n815 ^ n809 ;
  assign n821 = n817 ^ n806 ;
  assign n988 = n987 ^ n821 ;
  assign n508 = n487 ^ n483 ;
  assign n509 = n488 ^ n484 ;
  assign n511 = n508 & n509 ;
  assign n506 = n485 ^ n481 ;
  assign n507 = n486 ^ n482 ;
  assign n510 = n506 & n507 ;
  assign n515 = n511 ^ n510 ;
  assign n520 = n518 ^ n515 ;
  assign n521 = n520 ^ n504 ;
  assign n532 = n526 ^ n521 ;
  assign n479 = n477 ^ n472 ;
  assign n533 = n532 ^ n479 ;
  assign n556 = n542 ^ n533 ;
  assign n386 = n384 ^ n378 ;
  assign n390 = n386 ^ n375 ;
  assign n557 = n556 ^ n390 ;
  assign n1483 = n988 ^ n557 ;
  assign n4402 = n2871 ^ n1483 ;
  assign n2331 = n2327 ^ n2325 ;
  assign n2332 = n2328 ^ n2326 ;
  assign n2333 = n2331 & n2332 ;
  assign n2335 = n2334 ^ n2333 ;
  assign n2336 = n2335 ^ n2330 ;
  assign n2341 = n2338 ^ n2336 ;
  assign n2324 = n2323 ^ n2321 ;
  assign n2342 = n2341 ^ n2324 ;
  assign n2353 = n2346 ^ n2342 ;
  assign n2297 = n2296 ^ n2294 ;
  assign n2299 = n2297 ^ n2292 ;
  assign n2354 = n2353 ^ n2299 ;
  assign n2377 = n2362 ^ n2354 ;
  assign n2204 = n2203 ^ n2201 ;
  assign n2206 = n2204 ^ n2199 ;
  assign n2210 = n2206 ^ n2195 ;
  assign n2378 = n2377 ^ n2210 ;
  assign n1900 = n1896 ^ n1894 ;
  assign n1901 = n1897 ^ n1895 ;
  assign n1902 = n1900 & n1901 ;
  assign n1904 = n1903 ^ n1902 ;
  assign n1905 = n1904 ^ n1899 ;
  assign n1910 = n1907 ^ n1905 ;
  assign n1893 = n1892 ^ n1890 ;
  assign n1911 = n1910 ^ n1893 ;
  assign n1922 = n1915 ^ n1911 ;
  assign n1866 = n1865 ^ n1863 ;
  assign n1868 = n1866 ^ n1861 ;
  assign n1923 = n1922 ^ n1868 ;
  assign n1946 = n1931 ^ n1923 ;
  assign n1773 = n1772 ^ n1770 ;
  assign n1775 = n1773 ^ n1768 ;
  assign n1779 = n1775 ^ n1764 ;
  assign n1947 = n1946 ^ n1779 ;
  assign n2872 = n2378 ^ n1947 ;
  assign n943 = n939 ^ n937 ;
  assign n944 = n940 ^ n938 ;
  assign n945 = n943 & n944 ;
  assign n947 = n946 ^ n945 ;
  assign n948 = n947 ^ n942 ;
  assign n953 = n950 ^ n948 ;
  assign n936 = n935 ^ n933 ;
  assign n954 = n953 ^ n936 ;
  assign n965 = n958 ^ n954 ;
  assign n909 = n908 ^ n906 ;
  assign n911 = n909 ^ n904 ;
  assign n966 = n965 ^ n911 ;
  assign n989 = n974 ^ n966 ;
  assign n816 = n815 ^ n813 ;
  assign n818 = n816 ^ n811 ;
  assign n822 = n818 ^ n807 ;
  assign n990 = n989 ^ n822 ;
  assign n512 = n508 ^ n506 ;
  assign n513 = n509 ^ n507 ;
  assign n514 = n512 & n513 ;
  assign n516 = n515 ^ n514 ;
  assign n517 = n516 ^ n511 ;
  assign n522 = n519 ^ n517 ;
  assign n505 = n504 ^ n502 ;
  assign n523 = n522 ^ n505 ;
  assign n534 = n527 ^ n523 ;
  assign n478 = n477 ^ n475 ;
  assign n480 = n478 ^ n473 ;
  assign n535 = n534 ^ n480 ;
  assign n558 = n543 ^ n535 ;
  assign n385 = n384 ^ n382 ;
  assign n387 = n385 ^ n380 ;
  assign n391 = n387 ^ n376 ;
  assign n559 = n558 ^ n391 ;
  assign n1484 = n990 ^ n559 ;
  assign n4403 = n2872 ^ n1484 ;
  assign n2424 = x63 ^ x47 ;
  assign n2425 = x127 ^ x111 ;
  assign n2598 = n2424 & n2425 ;
  assign n2422 = x62 ^ x46 ;
  assign n2423 = x126 ^ x110 ;
  assign n2597 = n2422 & n2423 ;
  assign n2602 = n2598 ^ n2597 ;
  assign n2420 = x61 ^ x45 ;
  assign n2421 = x125 ^ x109 ;
  assign n2590 = n2420 & n2421 ;
  assign n2418 = x60 ^ x44 ;
  assign n2419 = x124 ^ x108 ;
  assign n2589 = n2418 & n2419 ;
  assign n2594 = n2590 ^ n2589 ;
  assign n2618 = n2602 ^ n2594 ;
  assign n2416 = x59 ^ x43 ;
  assign n2417 = x123 ^ x107 ;
  assign n2563 = n2416 & n2417 ;
  assign n2414 = x58 ^ x42 ;
  assign n2415 = x122 ^ x106 ;
  assign n2562 = n2414 & n2415 ;
  assign n2567 = n2563 ^ n2562 ;
  assign n2412 = x57 ^ x41 ;
  assign n2413 = x121 ^ x105 ;
  assign n2555 = n2412 & n2413 ;
  assign n2410 = x56 ^ x40 ;
  assign n2411 = x120 ^ x104 ;
  assign n2554 = n2410 & n2411 ;
  assign n2559 = n2555 ^ n2554 ;
  assign n2583 = n2567 ^ n2559 ;
  assign n2670 = n2618 ^ n2583 ;
  assign n2408 = x55 ^ x39 ;
  assign n2409 = x119 ^ x103 ;
  assign n2470 = n2408 & n2409 ;
  assign n2406 = x54 ^ x38 ;
  assign n2407 = x118 ^ x102 ;
  assign n2469 = n2406 & n2407 ;
  assign n2474 = n2470 ^ n2469 ;
  assign n2404 = x53 ^ x37 ;
  assign n2405 = x117 ^ x101 ;
  assign n2462 = n2404 & n2405 ;
  assign n2402 = x52 ^ x36 ;
  assign n2403 = x116 ^ x100 ;
  assign n2461 = n2402 & n2403 ;
  assign n2466 = n2462 ^ n2461 ;
  assign n2490 = n2474 ^ n2466 ;
  assign n2400 = x51 ^ x35 ;
  assign n2401 = x115 ^ x99 ;
  assign n2435 = n2400 & n2401 ;
  assign n2398 = x50 ^ x34 ;
  assign n2399 = x114 ^ x98 ;
  assign n2434 = n2398 & n2399 ;
  assign n2439 = n2435 ^ n2434 ;
  assign n2396 = x49 ^ x33 ;
  assign n2397 = x113 ^ x97 ;
  assign n2427 = n2396 & n2397 ;
  assign n2394 = x48 ^ x32 ;
  assign n2395 = x112 ^ x96 ;
  assign n2426 = n2394 & n2395 ;
  assign n2431 = n2427 ^ n2426 ;
  assign n2455 = n2439 ^ n2431 ;
  assign n2542 = n2490 ^ n2455 ;
  assign n2833 = n2670 ^ n2542 ;
  assign n2873 = n2857 ^ n2833 ;
  assign n2874 = n2873 ^ n2364 ;
  assign n1036 = x31 ^ x15 ;
  assign n1037 = x95 ^ x79 ;
  assign n1210 = n1036 & n1037 ;
  assign n1034 = x30 ^ x14 ;
  assign n1035 = x94 ^ x78 ;
  assign n1209 = n1034 & n1035 ;
  assign n1214 = n1210 ^ n1209 ;
  assign n1032 = x29 ^ x13 ;
  assign n1033 = x93 ^ x77 ;
  assign n1202 = n1032 & n1033 ;
  assign n1030 = x28 ^ x12 ;
  assign n1031 = x92 ^ x76 ;
  assign n1201 = n1030 & n1031 ;
  assign n1206 = n1202 ^ n1201 ;
  assign n1230 = n1214 ^ n1206 ;
  assign n1028 = x27 ^ x11 ;
  assign n1029 = x91 ^ x75 ;
  assign n1175 = n1028 & n1029 ;
  assign n1026 = x26 ^ x10 ;
  assign n1027 = x90 ^ x74 ;
  assign n1174 = n1026 & n1027 ;
  assign n1179 = n1175 ^ n1174 ;
  assign n1024 = x25 ^ x9 ;
  assign n1025 = x89 ^ x73 ;
  assign n1167 = n1024 & n1025 ;
  assign n1022 = x24 ^ x8 ;
  assign n1023 = x88 ^ x72 ;
  assign n1166 = n1022 & n1023 ;
  assign n1171 = n1167 ^ n1166 ;
  assign n1195 = n1179 ^ n1171 ;
  assign n1282 = n1230 ^ n1195 ;
  assign n1020 = x23 ^ x7 ;
  assign n1021 = x87 ^ x71 ;
  assign n1082 = n1020 & n1021 ;
  assign n1018 = x22 ^ x6 ;
  assign n1019 = x86 ^ x70 ;
  assign n1081 = n1018 & n1019 ;
  assign n1086 = n1082 ^ n1081 ;
  assign n1016 = x21 ^ x5 ;
  assign n1017 = x85 ^ x69 ;
  assign n1074 = n1016 & n1017 ;
  assign n1014 = x20 ^ x4 ;
  assign n1015 = x84 ^ x68 ;
  assign n1073 = n1014 & n1015 ;
  assign n1078 = n1074 ^ n1073 ;
  assign n1102 = n1086 ^ n1078 ;
  assign n1012 = x19 ^ x3 ;
  assign n1013 = x83 ^ x67 ;
  assign n1047 = n1012 & n1013 ;
  assign n1010 = x18 ^ x2 ;
  assign n1011 = x82 ^ x66 ;
  assign n1046 = n1010 & n1011 ;
  assign n1051 = n1047 ^ n1046 ;
  assign n1008 = x17 ^ x1 ;
  assign n1009 = x81 ^ x65 ;
  assign n1039 = n1008 & n1009 ;
  assign n1006 = x16 ^ x0 ;
  assign n1007 = x80 ^ x64 ;
  assign n1038 = n1006 & n1007 ;
  assign n1043 = n1039 ^ n1038 ;
  assign n1067 = n1051 ^ n1043 ;
  assign n1154 = n1102 ^ n1067 ;
  assign n1445 = n1282 ^ n1154 ;
  assign n1485 = n1469 ^ n1445 ;
  assign n1486 = n1485 ^ n976 ;
  assign n4404 = n2874 ^ n1486 ;
  assign n2599 = n2424 ^ n2422 ;
  assign n2600 = n2425 ^ n2423 ;
  assign n2601 = n2599 & n2600 ;
  assign n2603 = n2602 ^ n2601 ;
  assign n2604 = n2603 ^ n2598 ;
  assign n2591 = n2420 ^ n2418 ;
  assign n2592 = n2421 ^ n2419 ;
  assign n2593 = n2591 & n2592 ;
  assign n2595 = n2594 ^ n2593 ;
  assign n2596 = n2595 ^ n2590 ;
  assign n2619 = n2604 ^ n2596 ;
  assign n2564 = n2416 ^ n2414 ;
  assign n2565 = n2417 ^ n2415 ;
  assign n2566 = n2564 & n2565 ;
  assign n2568 = n2567 ^ n2566 ;
  assign n2569 = n2568 ^ n2563 ;
  assign n2556 = n2412 ^ n2410 ;
  assign n2557 = n2413 ^ n2411 ;
  assign n2558 = n2556 & n2557 ;
  assign n2560 = n2559 ^ n2558 ;
  assign n2561 = n2560 ^ n2555 ;
  assign n2584 = n2569 ^ n2561 ;
  assign n2671 = n2619 ^ n2584 ;
  assign n2471 = n2408 ^ n2406 ;
  assign n2472 = n2409 ^ n2407 ;
  assign n2473 = n2471 & n2472 ;
  assign n2475 = n2474 ^ n2473 ;
  assign n2476 = n2475 ^ n2470 ;
  assign n2463 = n2404 ^ n2402 ;
  assign n2464 = n2405 ^ n2403 ;
  assign n2465 = n2463 & n2464 ;
  assign n2467 = n2466 ^ n2465 ;
  assign n2468 = n2467 ^ n2462 ;
  assign n2491 = n2476 ^ n2468 ;
  assign n2436 = n2400 ^ n2398 ;
  assign n2437 = n2401 ^ n2399 ;
  assign n2438 = n2436 & n2437 ;
  assign n2440 = n2439 ^ n2438 ;
  assign n2441 = n2440 ^ n2435 ;
  assign n2428 = n2396 ^ n2394 ;
  assign n2429 = n2397 ^ n2395 ;
  assign n2430 = n2428 & n2429 ;
  assign n2432 = n2431 ^ n2430 ;
  assign n2433 = n2432 ^ n2427 ;
  assign n2456 = n2441 ^ n2433 ;
  assign n2543 = n2491 ^ n2456 ;
  assign n2834 = n2671 ^ n2543 ;
  assign n2875 = n2858 ^ n2834 ;
  assign n2876 = n2875 ^ n2366 ;
  assign n1211 = n1036 ^ n1034 ;
  assign n1212 = n1037 ^ n1035 ;
  assign n1213 = n1211 & n1212 ;
  assign n1215 = n1214 ^ n1213 ;
  assign n1216 = n1215 ^ n1210 ;
  assign n1203 = n1032 ^ n1030 ;
  assign n1204 = n1033 ^ n1031 ;
  assign n1205 = n1203 & n1204 ;
  assign n1207 = n1206 ^ n1205 ;
  assign n1208 = n1207 ^ n1202 ;
  assign n1231 = n1216 ^ n1208 ;
  assign n1176 = n1028 ^ n1026 ;
  assign n1177 = n1029 ^ n1027 ;
  assign n1178 = n1176 & n1177 ;
  assign n1180 = n1179 ^ n1178 ;
  assign n1181 = n1180 ^ n1175 ;
  assign n1168 = n1024 ^ n1022 ;
  assign n1169 = n1025 ^ n1023 ;
  assign n1170 = n1168 & n1169 ;
  assign n1172 = n1171 ^ n1170 ;
  assign n1173 = n1172 ^ n1167 ;
  assign n1196 = n1181 ^ n1173 ;
  assign n1283 = n1231 ^ n1196 ;
  assign n1083 = n1020 ^ n1018 ;
  assign n1084 = n1021 ^ n1019 ;
  assign n1085 = n1083 & n1084 ;
  assign n1087 = n1086 ^ n1085 ;
  assign n1088 = n1087 ^ n1082 ;
  assign n1075 = n1016 ^ n1014 ;
  assign n1076 = n1017 ^ n1015 ;
  assign n1077 = n1075 & n1076 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n1080 = n1079 ^ n1074 ;
  assign n1103 = n1088 ^ n1080 ;
  assign n1048 = n1012 ^ n1010 ;
  assign n1049 = n1013 ^ n1011 ;
  assign n1050 = n1048 & n1049 ;
  assign n1052 = n1051 ^ n1050 ;
  assign n1053 = n1052 ^ n1047 ;
  assign n1040 = n1008 ^ n1006 ;
  assign n1041 = n1009 ^ n1007 ;
  assign n1042 = n1040 & n1041 ;
  assign n1044 = n1043 ^ n1042 ;
  assign n1045 = n1044 ^ n1039 ;
  assign n1068 = n1053 ^ n1045 ;
  assign n1155 = n1103 ^ n1068 ;
  assign n1446 = n1283 ^ n1155 ;
  assign n1487 = n1470 ^ n1446 ;
  assign n1488 = n1487 ^ n978 ;
  assign n4405 = n2876 ^ n1488 ;
  assign n2608 = n2424 ^ n2420 ;
  assign n2609 = n2425 ^ n2421 ;
  assign n2611 = n2608 & n2609 ;
  assign n2606 = n2422 ^ n2418 ;
  assign n2607 = n2423 ^ n2419 ;
  assign n2610 = n2606 & n2607 ;
  assign n2615 = n2611 ^ n2610 ;
  assign n2620 = n2618 ^ n2615 ;
  assign n2621 = n2620 ^ n2604 ;
  assign n2573 = n2416 ^ n2412 ;
  assign n2574 = n2417 ^ n2413 ;
  assign n2576 = n2573 & n2574 ;
  assign n2571 = n2414 ^ n2410 ;
  assign n2572 = n2415 ^ n2411 ;
  assign n2575 = n2571 & n2572 ;
  assign n2580 = n2576 ^ n2575 ;
  assign n2585 = n2583 ^ n2580 ;
  assign n2586 = n2585 ^ n2569 ;
  assign n2672 = n2621 ^ n2586 ;
  assign n2480 = n2408 ^ n2404 ;
  assign n2481 = n2409 ^ n2405 ;
  assign n2483 = n2480 & n2481 ;
  assign n2478 = n2406 ^ n2402 ;
  assign n2479 = n2407 ^ n2403 ;
  assign n2482 = n2478 & n2479 ;
  assign n2487 = n2483 ^ n2482 ;
  assign n2492 = n2490 ^ n2487 ;
  assign n2493 = n2492 ^ n2476 ;
  assign n2445 = n2400 ^ n2396 ;
  assign n2446 = n2401 ^ n2397 ;
  assign n2448 = n2445 & n2446 ;
  assign n2443 = n2398 ^ n2394 ;
  assign n2444 = n2399 ^ n2395 ;
  assign n2447 = n2443 & n2444 ;
  assign n2452 = n2448 ^ n2447 ;
  assign n2457 = n2455 ^ n2452 ;
  assign n2458 = n2457 ^ n2441 ;
  assign n2544 = n2493 ^ n2458 ;
  assign n2835 = n2672 ^ n2544 ;
  assign n2877 = n2859 ^ n2835 ;
  assign n2878 = n2877 ^ n2368 ;
  assign n1220 = n1036 ^ n1032 ;
  assign n1221 = n1037 ^ n1033 ;
  assign n1223 = n1220 & n1221 ;
  assign n1218 = n1034 ^ n1030 ;
  assign n1219 = n1035 ^ n1031 ;
  assign n1222 = n1218 & n1219 ;
  assign n1227 = n1223 ^ n1222 ;
  assign n1232 = n1230 ^ n1227 ;
  assign n1233 = n1232 ^ n1216 ;
  assign n1185 = n1028 ^ n1024 ;
  assign n1186 = n1029 ^ n1025 ;
  assign n1188 = n1185 & n1186 ;
  assign n1183 = n1026 ^ n1022 ;
  assign n1184 = n1027 ^ n1023 ;
  assign n1187 = n1183 & n1184 ;
  assign n1192 = n1188 ^ n1187 ;
  assign n1197 = n1195 ^ n1192 ;
  assign n1198 = n1197 ^ n1181 ;
  assign n1284 = n1233 ^ n1198 ;
  assign n1092 = n1020 ^ n1016 ;
  assign n1093 = n1021 ^ n1017 ;
  assign n1095 = n1092 & n1093 ;
  assign n1090 = n1018 ^ n1014 ;
  assign n1091 = n1019 ^ n1015 ;
  assign n1094 = n1090 & n1091 ;
  assign n1099 = n1095 ^ n1094 ;
  assign n1104 = n1102 ^ n1099 ;
  assign n1105 = n1104 ^ n1088 ;
  assign n1057 = n1012 ^ n1008 ;
  assign n1058 = n1013 ^ n1009 ;
  assign n1060 = n1057 & n1058 ;
  assign n1055 = n1010 ^ n1006 ;
  assign n1056 = n1011 ^ n1007 ;
  assign n1059 = n1055 & n1056 ;
  assign n1064 = n1060 ^ n1059 ;
  assign n1069 = n1067 ^ n1064 ;
  assign n1070 = n1069 ^ n1053 ;
  assign n1156 = n1105 ^ n1070 ;
  assign n1447 = n1284 ^ n1156 ;
  assign n1489 = n1471 ^ n1447 ;
  assign n1490 = n1489 ^ n980 ;
  assign n4406 = n2878 ^ n1490 ;
  assign n2612 = n2608 ^ n2606 ;
  assign n2613 = n2609 ^ n2607 ;
  assign n2614 = n2612 & n2613 ;
  assign n2616 = n2615 ^ n2614 ;
  assign n2617 = n2616 ^ n2611 ;
  assign n2622 = n2619 ^ n2617 ;
  assign n2605 = n2604 ^ n2602 ;
  assign n2623 = n2622 ^ n2605 ;
  assign n2577 = n2573 ^ n2571 ;
  assign n2578 = n2574 ^ n2572 ;
  assign n2579 = n2577 & n2578 ;
  assign n2581 = n2580 ^ n2579 ;
  assign n2582 = n2581 ^ n2576 ;
  assign n2587 = n2584 ^ n2582 ;
  assign n2570 = n2569 ^ n2567 ;
  assign n2588 = n2587 ^ n2570 ;
  assign n2673 = n2623 ^ n2588 ;
  assign n2484 = n2480 ^ n2478 ;
  assign n2485 = n2481 ^ n2479 ;
  assign n2486 = n2484 & n2485 ;
  assign n2488 = n2487 ^ n2486 ;
  assign n2489 = n2488 ^ n2483 ;
  assign n2494 = n2491 ^ n2489 ;
  assign n2477 = n2476 ^ n2474 ;
  assign n2495 = n2494 ^ n2477 ;
  assign n2449 = n2445 ^ n2443 ;
  assign n2450 = n2446 ^ n2444 ;
  assign n2451 = n2449 & n2450 ;
  assign n2453 = n2452 ^ n2451 ;
  assign n2454 = n2453 ^ n2448 ;
  assign n2459 = n2456 ^ n2454 ;
  assign n2442 = n2441 ^ n2439 ;
  assign n2460 = n2459 ^ n2442 ;
  assign n2545 = n2495 ^ n2460 ;
  assign n2836 = n2673 ^ n2545 ;
  assign n2879 = n2860 ^ n2836 ;
  assign n2880 = n2879 ^ n2370 ;
  assign n1224 = n1220 ^ n1218 ;
  assign n1225 = n1221 ^ n1219 ;
  assign n1226 = n1224 & n1225 ;
  assign n1228 = n1227 ^ n1226 ;
  assign n1229 = n1228 ^ n1223 ;
  assign n1234 = n1231 ^ n1229 ;
  assign n1217 = n1216 ^ n1214 ;
  assign n1235 = n1234 ^ n1217 ;
  assign n1189 = n1185 ^ n1183 ;
  assign n1190 = n1186 ^ n1184 ;
  assign n1191 = n1189 & n1190 ;
  assign n1193 = n1192 ^ n1191 ;
  assign n1194 = n1193 ^ n1188 ;
  assign n1199 = n1196 ^ n1194 ;
  assign n1182 = n1181 ^ n1179 ;
  assign n1200 = n1199 ^ n1182 ;
  assign n1285 = n1235 ^ n1200 ;
  assign n1096 = n1092 ^ n1090 ;
  assign n1097 = n1093 ^ n1091 ;
  assign n1098 = n1096 & n1097 ;
  assign n1100 = n1099 ^ n1098 ;
  assign n1101 = n1100 ^ n1095 ;
  assign n1106 = n1103 ^ n1101 ;
  assign n1089 = n1088 ^ n1086 ;
  assign n1107 = n1106 ^ n1089 ;
  assign n1061 = n1057 ^ n1055 ;
  assign n1062 = n1058 ^ n1056 ;
  assign n1063 = n1061 & n1062 ;
  assign n1065 = n1064 ^ n1063 ;
  assign n1066 = n1065 ^ n1060 ;
  assign n1071 = n1068 ^ n1066 ;
  assign n1054 = n1053 ^ n1051 ;
  assign n1072 = n1071 ^ n1054 ;
  assign n1157 = n1107 ^ n1072 ;
  assign n1448 = n1285 ^ n1157 ;
  assign n1491 = n1472 ^ n1448 ;
  assign n1492 = n1491 ^ n982 ;
  assign n4407 = n2880 ^ n1492 ;
  assign n2633 = n2424 ^ n2416 ;
  assign n2634 = n2425 ^ n2417 ;
  assign n2644 = n2633 & n2634 ;
  assign n2631 = n2422 ^ n2414 ;
  assign n2632 = n2423 ^ n2415 ;
  assign n2643 = n2631 & n2632 ;
  assign n2648 = n2644 ^ n2643 ;
  assign n2629 = n2420 ^ n2412 ;
  assign n2630 = n2421 ^ n2413 ;
  assign n2636 = n2629 & n2630 ;
  assign n2627 = n2418 ^ n2410 ;
  assign n2628 = n2419 ^ n2411 ;
  assign n2635 = n2627 & n2628 ;
  assign n2640 = n2636 ^ n2635 ;
  assign n2664 = n2648 ^ n2640 ;
  assign n2674 = n2670 ^ n2664 ;
  assign n2675 = n2674 ^ n2621 ;
  assign n2505 = n2408 ^ n2400 ;
  assign n2506 = n2409 ^ n2401 ;
  assign n2516 = n2505 & n2506 ;
  assign n2503 = n2406 ^ n2398 ;
  assign n2504 = n2407 ^ n2399 ;
  assign n2515 = n2503 & n2504 ;
  assign n2520 = n2516 ^ n2515 ;
  assign n2501 = n2404 ^ n2396 ;
  assign n2502 = n2405 ^ n2397 ;
  assign n2508 = n2501 & n2502 ;
  assign n2499 = n2402 ^ n2394 ;
  assign n2500 = n2403 ^ n2395 ;
  assign n2507 = n2499 & n2500 ;
  assign n2512 = n2508 ^ n2507 ;
  assign n2536 = n2520 ^ n2512 ;
  assign n2546 = n2542 ^ n2536 ;
  assign n2547 = n2546 ^ n2493 ;
  assign n2837 = n2675 ^ n2547 ;
  assign n2881 = n2861 ^ n2837 ;
  assign n2882 = n2881 ^ n2372 ;
  assign n1245 = n1036 ^ n1028 ;
  assign n1246 = n1037 ^ n1029 ;
  assign n1256 = n1245 & n1246 ;
  assign n1243 = n1034 ^ n1026 ;
  assign n1244 = n1035 ^ n1027 ;
  assign n1255 = n1243 & n1244 ;
  assign n1260 = n1256 ^ n1255 ;
  assign n1241 = n1032 ^ n1024 ;
  assign n1242 = n1033 ^ n1025 ;
  assign n1248 = n1241 & n1242 ;
  assign n1239 = n1030 ^ n1022 ;
  assign n1240 = n1031 ^ n1023 ;
  assign n1247 = n1239 & n1240 ;
  assign n1252 = n1248 ^ n1247 ;
  assign n1276 = n1260 ^ n1252 ;
  assign n1286 = n1282 ^ n1276 ;
  assign n1287 = n1286 ^ n1233 ;
  assign n1117 = n1020 ^ n1012 ;
  assign n1118 = n1021 ^ n1013 ;
  assign n1128 = n1117 & n1118 ;
  assign n1115 = n1018 ^ n1010 ;
  assign n1116 = n1019 ^ n1011 ;
  assign n1127 = n1115 & n1116 ;
  assign n1132 = n1128 ^ n1127 ;
  assign n1113 = n1016 ^ n1008 ;
  assign n1114 = n1017 ^ n1009 ;
  assign n1120 = n1113 & n1114 ;
  assign n1111 = n1014 ^ n1006 ;
  assign n1112 = n1015 ^ n1007 ;
  assign n1119 = n1111 & n1112 ;
  assign n1124 = n1120 ^ n1119 ;
  assign n1148 = n1132 ^ n1124 ;
  assign n1158 = n1154 ^ n1148 ;
  assign n1159 = n1158 ^ n1105 ;
  assign n1449 = n1287 ^ n1159 ;
  assign n1493 = n1473 ^ n1449 ;
  assign n1494 = n1493 ^ n984 ;
  assign n4408 = n2882 ^ n1494 ;
  assign n2645 = n2633 ^ n2631 ;
  assign n2646 = n2634 ^ n2632 ;
  assign n2647 = n2645 & n2646 ;
  assign n2649 = n2648 ^ n2647 ;
  assign n2650 = n2649 ^ n2644 ;
  assign n2637 = n2629 ^ n2627 ;
  assign n2638 = n2630 ^ n2628 ;
  assign n2639 = n2637 & n2638 ;
  assign n2641 = n2640 ^ n2639 ;
  assign n2642 = n2641 ^ n2636 ;
  assign n2665 = n2650 ^ n2642 ;
  assign n2676 = n2671 ^ n2665 ;
  assign n2677 = n2676 ^ n2623 ;
  assign n2517 = n2505 ^ n2503 ;
  assign n2518 = n2506 ^ n2504 ;
  assign n2519 = n2517 & n2518 ;
  assign n2521 = n2520 ^ n2519 ;
  assign n2522 = n2521 ^ n2516 ;
  assign n2509 = n2501 ^ n2499 ;
  assign n2510 = n2502 ^ n2500 ;
  assign n2511 = n2509 & n2510 ;
  assign n2513 = n2512 ^ n2511 ;
  assign n2514 = n2513 ^ n2508 ;
  assign n2537 = n2522 ^ n2514 ;
  assign n2548 = n2543 ^ n2537 ;
  assign n2549 = n2548 ^ n2495 ;
  assign n2838 = n2677 ^ n2549 ;
  assign n2883 = n2862 ^ n2838 ;
  assign n2884 = n2883 ^ n2374 ;
  assign n1257 = n1245 ^ n1243 ;
  assign n1258 = n1246 ^ n1244 ;
  assign n1259 = n1257 & n1258 ;
  assign n1261 = n1260 ^ n1259 ;
  assign n1262 = n1261 ^ n1256 ;
  assign n1249 = n1241 ^ n1239 ;
  assign n1250 = n1242 ^ n1240 ;
  assign n1251 = n1249 & n1250 ;
  assign n1253 = n1252 ^ n1251 ;
  assign n1254 = n1253 ^ n1248 ;
  assign n1277 = n1262 ^ n1254 ;
  assign n1288 = n1283 ^ n1277 ;
  assign n1289 = n1288 ^ n1235 ;
  assign n1129 = n1117 ^ n1115 ;
  assign n1130 = n1118 ^ n1116 ;
  assign n1131 = n1129 & n1130 ;
  assign n1133 = n1132 ^ n1131 ;
  assign n1134 = n1133 ^ n1128 ;
  assign n1121 = n1113 ^ n1111 ;
  assign n1122 = n1114 ^ n1112 ;
  assign n1123 = n1121 & n1122 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1126 = n1125 ^ n1120 ;
  assign n1149 = n1134 ^ n1126 ;
  assign n1160 = n1155 ^ n1149 ;
  assign n1161 = n1160 ^ n1107 ;
  assign n1450 = n1289 ^ n1161 ;
  assign n1495 = n1474 ^ n1450 ;
  assign n1496 = n1495 ^ n986 ;
  assign n4409 = n2884 ^ n1496 ;
  assign n2654 = n2633 ^ n2629 ;
  assign n2655 = n2634 ^ n2630 ;
  assign n2657 = n2654 & n2655 ;
  assign n2652 = n2631 ^ n2627 ;
  assign n2653 = n2632 ^ n2628 ;
  assign n2656 = n2652 & n2653 ;
  assign n2661 = n2657 ^ n2656 ;
  assign n2666 = n2664 ^ n2661 ;
  assign n2667 = n2666 ^ n2650 ;
  assign n2678 = n2672 ^ n2667 ;
  assign n2625 = n2623 ^ n2618 ;
  assign n2679 = n2678 ^ n2625 ;
  assign n2526 = n2505 ^ n2501 ;
  assign n2527 = n2506 ^ n2502 ;
  assign n2529 = n2526 & n2527 ;
  assign n2524 = n2503 ^ n2499 ;
  assign n2525 = n2504 ^ n2500 ;
  assign n2528 = n2524 & n2525 ;
  assign n2533 = n2529 ^ n2528 ;
  assign n2538 = n2536 ^ n2533 ;
  assign n2539 = n2538 ^ n2522 ;
  assign n2550 = n2544 ^ n2539 ;
  assign n2497 = n2495 ^ n2490 ;
  assign n2551 = n2550 ^ n2497 ;
  assign n2839 = n2679 ^ n2551 ;
  assign n2885 = n2863 ^ n2839 ;
  assign n2886 = n2885 ^ n2376 ;
  assign n1266 = n1245 ^ n1241 ;
  assign n1267 = n1246 ^ n1242 ;
  assign n1269 = n1266 & n1267 ;
  assign n1264 = n1243 ^ n1239 ;
  assign n1265 = n1244 ^ n1240 ;
  assign n1268 = n1264 & n1265 ;
  assign n1273 = n1269 ^ n1268 ;
  assign n1278 = n1276 ^ n1273 ;
  assign n1279 = n1278 ^ n1262 ;
  assign n1290 = n1284 ^ n1279 ;
  assign n1237 = n1235 ^ n1230 ;
  assign n1291 = n1290 ^ n1237 ;
  assign n1138 = n1117 ^ n1113 ;
  assign n1139 = n1118 ^ n1114 ;
  assign n1141 = n1138 & n1139 ;
  assign n1136 = n1115 ^ n1111 ;
  assign n1137 = n1116 ^ n1112 ;
  assign n1140 = n1136 & n1137 ;
  assign n1145 = n1141 ^ n1140 ;
  assign n1150 = n1148 ^ n1145 ;
  assign n1151 = n1150 ^ n1134 ;
  assign n1162 = n1156 ^ n1151 ;
  assign n1109 = n1107 ^ n1102 ;
  assign n1163 = n1162 ^ n1109 ;
  assign n1451 = n1291 ^ n1163 ;
  assign n1497 = n1475 ^ n1451 ;
  assign n1498 = n1497 ^ n988 ;
  assign n4410 = n2886 ^ n1498 ;
  assign n2658 = n2654 ^ n2652 ;
  assign n2659 = n2655 ^ n2653 ;
  assign n2660 = n2658 & n2659 ;
  assign n2662 = n2661 ^ n2660 ;
  assign n2663 = n2662 ^ n2657 ;
  assign n2668 = n2665 ^ n2663 ;
  assign n2651 = n2650 ^ n2648 ;
  assign n2669 = n2668 ^ n2651 ;
  assign n2680 = n2673 ^ n2669 ;
  assign n2624 = n2623 ^ n2621 ;
  assign n2626 = n2624 ^ n2619 ;
  assign n2681 = n2680 ^ n2626 ;
  assign n2530 = n2526 ^ n2524 ;
  assign n2531 = n2527 ^ n2525 ;
  assign n2532 = n2530 & n2531 ;
  assign n2534 = n2533 ^ n2532 ;
  assign n2535 = n2534 ^ n2529 ;
  assign n2540 = n2537 ^ n2535 ;
  assign n2523 = n2522 ^ n2520 ;
  assign n2541 = n2540 ^ n2523 ;
  assign n2552 = n2545 ^ n2541 ;
  assign n2496 = n2495 ^ n2493 ;
  assign n2498 = n2496 ^ n2491 ;
  assign n2553 = n2552 ^ n2498 ;
  assign n2840 = n2681 ^ n2553 ;
  assign n2887 = n2864 ^ n2840 ;
  assign n2888 = n2887 ^ n2378 ;
  assign n1270 = n1266 ^ n1264 ;
  assign n1271 = n1267 ^ n1265 ;
  assign n1272 = n1270 & n1271 ;
  assign n1274 = n1273 ^ n1272 ;
  assign n1275 = n1274 ^ n1269 ;
  assign n1280 = n1277 ^ n1275 ;
  assign n1263 = n1262 ^ n1260 ;
  assign n1281 = n1280 ^ n1263 ;
  assign n1292 = n1285 ^ n1281 ;
  assign n1236 = n1235 ^ n1233 ;
  assign n1238 = n1236 ^ n1231 ;
  assign n1293 = n1292 ^ n1238 ;
  assign n1142 = n1138 ^ n1136 ;
  assign n1143 = n1139 ^ n1137 ;
  assign n1144 = n1142 & n1143 ;
  assign n1146 = n1145 ^ n1144 ;
  assign n1147 = n1146 ^ n1141 ;
  assign n1152 = n1149 ^ n1147 ;
  assign n1135 = n1134 ^ n1132 ;
  assign n1153 = n1152 ^ n1135 ;
  assign n1164 = n1157 ^ n1153 ;
  assign n1108 = n1107 ^ n1105 ;
  assign n1110 = n1108 ^ n1103 ;
  assign n1165 = n1164 ^ n1110 ;
  assign n1452 = n1293 ^ n1165 ;
  assign n1499 = n1476 ^ n1452 ;
  assign n1500 = n1499 ^ n990 ;
  assign n4411 = n2888 ^ n1500 ;
  assign n2703 = n2424 ^ n2408 ;
  assign n2704 = n2425 ^ n2409 ;
  assign n2749 = n2703 & n2704 ;
  assign n2701 = n2422 ^ n2406 ;
  assign n2702 = n2423 ^ n2407 ;
  assign n2748 = n2701 & n2702 ;
  assign n2753 = n2749 ^ n2748 ;
  assign n2699 = n2420 ^ n2404 ;
  assign n2700 = n2421 ^ n2405 ;
  assign n2741 = n2699 & n2700 ;
  assign n2697 = n2418 ^ n2402 ;
  assign n2698 = n2419 ^ n2403 ;
  assign n2740 = n2697 & n2698 ;
  assign n2745 = n2741 ^ n2740 ;
  assign n2769 = n2753 ^ n2745 ;
  assign n2695 = n2416 ^ n2400 ;
  assign n2696 = n2417 ^ n2401 ;
  assign n2714 = n2695 & n2696 ;
  assign n2693 = n2414 ^ n2398 ;
  assign n2694 = n2415 ^ n2399 ;
  assign n2713 = n2693 & n2694 ;
  assign n2718 = n2714 ^ n2713 ;
  assign n2691 = n2412 ^ n2396 ;
  assign n2692 = n2413 ^ n2397 ;
  assign n2706 = n2691 & n2692 ;
  assign n2689 = n2410 ^ n2394 ;
  assign n2690 = n2411 ^ n2395 ;
  assign n2705 = n2689 & n2690 ;
  assign n2710 = n2706 ^ n2705 ;
  assign n2734 = n2718 ^ n2710 ;
  assign n2821 = n2769 ^ n2734 ;
  assign n2841 = n2833 ^ n2821 ;
  assign n2842 = n2841 ^ n2675 ;
  assign n2889 = n2865 ^ n2842 ;
  assign n2386 = n2372 ^ n2355 ;
  assign n2890 = n2889 ^ n2386 ;
  assign n1315 = n1036 ^ n1020 ;
  assign n1316 = n1037 ^ n1021 ;
  assign n1361 = n1315 & n1316 ;
  assign n1313 = n1034 ^ n1018 ;
  assign n1314 = n1035 ^ n1019 ;
  assign n1360 = n1313 & n1314 ;
  assign n1365 = n1361 ^ n1360 ;
  assign n1311 = n1032 ^ n1016 ;
  assign n1312 = n1033 ^ n1017 ;
  assign n1353 = n1311 & n1312 ;
  assign n1309 = n1030 ^ n1014 ;
  assign n1310 = n1031 ^ n1015 ;
  assign n1352 = n1309 & n1310 ;
  assign n1357 = n1353 ^ n1352 ;
  assign n1381 = n1365 ^ n1357 ;
  assign n1307 = n1028 ^ n1012 ;
  assign n1308 = n1029 ^ n1013 ;
  assign n1326 = n1307 & n1308 ;
  assign n1305 = n1026 ^ n1010 ;
  assign n1306 = n1027 ^ n1011 ;
  assign n1325 = n1305 & n1306 ;
  assign n1330 = n1326 ^ n1325 ;
  assign n1303 = n1024 ^ n1008 ;
  assign n1304 = n1025 ^ n1009 ;
  assign n1318 = n1303 & n1304 ;
  assign n1301 = n1022 ^ n1006 ;
  assign n1302 = n1023 ^ n1007 ;
  assign n1317 = n1301 & n1302 ;
  assign n1322 = n1318 ^ n1317 ;
  assign n1346 = n1330 ^ n1322 ;
  assign n1433 = n1381 ^ n1346 ;
  assign n1453 = n1445 ^ n1433 ;
  assign n1454 = n1453 ^ n1287 ;
  assign n1501 = n1477 ^ n1454 ;
  assign n998 = n984 ^ n967 ;
  assign n1502 = n1501 ^ n998 ;
  assign n4412 = n2890 ^ n1502 ;
  assign n2750 = n2703 ^ n2701 ;
  assign n2751 = n2704 ^ n2702 ;
  assign n2752 = n2750 & n2751 ;
  assign n2754 = n2753 ^ n2752 ;
  assign n2755 = n2754 ^ n2749 ;
  assign n2742 = n2699 ^ n2697 ;
  assign n2743 = n2700 ^ n2698 ;
  assign n2744 = n2742 & n2743 ;
  assign n2746 = n2745 ^ n2744 ;
  assign n2747 = n2746 ^ n2741 ;
  assign n2770 = n2755 ^ n2747 ;
  assign n2715 = n2695 ^ n2693 ;
  assign n2716 = n2696 ^ n2694 ;
  assign n2717 = n2715 & n2716 ;
  assign n2719 = n2718 ^ n2717 ;
  assign n2720 = n2719 ^ n2714 ;
  assign n2707 = n2691 ^ n2689 ;
  assign n2708 = n2692 ^ n2690 ;
  assign n2709 = n2707 & n2708 ;
  assign n2711 = n2710 ^ n2709 ;
  assign n2712 = n2711 ^ n2706 ;
  assign n2735 = n2720 ^ n2712 ;
  assign n2822 = n2770 ^ n2735 ;
  assign n2843 = n2834 ^ n2822 ;
  assign n2844 = n2843 ^ n2677 ;
  assign n2891 = n2866 ^ n2844 ;
  assign n2387 = n2374 ^ n2356 ;
  assign n2892 = n2891 ^ n2387 ;
  assign n1362 = n1315 ^ n1313 ;
  assign n1363 = n1316 ^ n1314 ;
  assign n1364 = n1362 & n1363 ;
  assign n1366 = n1365 ^ n1364 ;
  assign n1367 = n1366 ^ n1361 ;
  assign n1354 = n1311 ^ n1309 ;
  assign n1355 = n1312 ^ n1310 ;
  assign n1356 = n1354 & n1355 ;
  assign n1358 = n1357 ^ n1356 ;
  assign n1359 = n1358 ^ n1353 ;
  assign n1382 = n1367 ^ n1359 ;
  assign n1327 = n1307 ^ n1305 ;
  assign n1328 = n1308 ^ n1306 ;
  assign n1329 = n1327 & n1328 ;
  assign n1331 = n1330 ^ n1329 ;
  assign n1332 = n1331 ^ n1326 ;
  assign n1319 = n1303 ^ n1301 ;
  assign n1320 = n1304 ^ n1302 ;
  assign n1321 = n1319 & n1320 ;
  assign n1323 = n1322 ^ n1321 ;
  assign n1324 = n1323 ^ n1318 ;
  assign n1347 = n1332 ^ n1324 ;
  assign n1434 = n1382 ^ n1347 ;
  assign n1455 = n1446 ^ n1434 ;
  assign n1456 = n1455 ^ n1289 ;
  assign n1503 = n1478 ^ n1456 ;
  assign n999 = n986 ^ n968 ;
  assign n1504 = n1503 ^ n999 ;
  assign n4413 = n2892 ^ n1504 ;
  assign n2759 = n2703 ^ n2699 ;
  assign n2760 = n2704 ^ n2700 ;
  assign n2762 = n2759 & n2760 ;
  assign n2757 = n2701 ^ n2697 ;
  assign n2758 = n2702 ^ n2698 ;
  assign n2761 = n2757 & n2758 ;
  assign n2766 = n2762 ^ n2761 ;
  assign n2771 = n2769 ^ n2766 ;
  assign n2772 = n2771 ^ n2755 ;
  assign n2724 = n2695 ^ n2691 ;
  assign n2725 = n2696 ^ n2692 ;
  assign n2727 = n2724 & n2725 ;
  assign n2722 = n2693 ^ n2689 ;
  assign n2723 = n2694 ^ n2690 ;
  assign n2726 = n2722 & n2723 ;
  assign n2731 = n2727 ^ n2726 ;
  assign n2736 = n2734 ^ n2731 ;
  assign n2737 = n2736 ^ n2720 ;
  assign n2823 = n2772 ^ n2737 ;
  assign n2845 = n2835 ^ n2823 ;
  assign n2846 = n2845 ^ n2679 ;
  assign n2893 = n2867 ^ n2846 ;
  assign n2388 = n2376 ^ n2357 ;
  assign n2894 = n2893 ^ n2388 ;
  assign n1371 = n1315 ^ n1311 ;
  assign n1372 = n1316 ^ n1312 ;
  assign n1374 = n1371 & n1372 ;
  assign n1369 = n1313 ^ n1309 ;
  assign n1370 = n1314 ^ n1310 ;
  assign n1373 = n1369 & n1370 ;
  assign n1378 = n1374 ^ n1373 ;
  assign n1383 = n1381 ^ n1378 ;
  assign n1384 = n1383 ^ n1367 ;
  assign n1336 = n1307 ^ n1303 ;
  assign n1337 = n1308 ^ n1304 ;
  assign n1339 = n1336 & n1337 ;
  assign n1334 = n1305 ^ n1301 ;
  assign n1335 = n1306 ^ n1302 ;
  assign n1338 = n1334 & n1335 ;
  assign n1343 = n1339 ^ n1338 ;
  assign n1348 = n1346 ^ n1343 ;
  assign n1349 = n1348 ^ n1332 ;
  assign n1435 = n1384 ^ n1349 ;
  assign n1457 = n1447 ^ n1435 ;
  assign n1458 = n1457 ^ n1291 ;
  assign n1505 = n1479 ^ n1458 ;
  assign n1000 = n988 ^ n969 ;
  assign n1506 = n1505 ^ n1000 ;
  assign n4414 = n2894 ^ n1506 ;
  assign n2763 = n2759 ^ n2757 ;
  assign n2764 = n2760 ^ n2758 ;
  assign n2765 = n2763 & n2764 ;
  assign n2767 = n2766 ^ n2765 ;
  assign n2768 = n2767 ^ n2762 ;
  assign n2773 = n2770 ^ n2768 ;
  assign n2756 = n2755 ^ n2753 ;
  assign n2774 = n2773 ^ n2756 ;
  assign n2728 = n2724 ^ n2722 ;
  assign n2729 = n2725 ^ n2723 ;
  assign n2730 = n2728 & n2729 ;
  assign n2732 = n2731 ^ n2730 ;
  assign n2733 = n2732 ^ n2727 ;
  assign n2738 = n2735 ^ n2733 ;
  assign n2721 = n2720 ^ n2718 ;
  assign n2739 = n2738 ^ n2721 ;
  assign n2824 = n2774 ^ n2739 ;
  assign n2847 = n2836 ^ n2824 ;
  assign n2848 = n2847 ^ n2681 ;
  assign n2895 = n2868 ^ n2848 ;
  assign n2389 = n2378 ^ n2358 ;
  assign n2896 = n2895 ^ n2389 ;
  assign n1375 = n1371 ^ n1369 ;
  assign n1376 = n1372 ^ n1370 ;
  assign n1377 = n1375 & n1376 ;
  assign n1379 = n1378 ^ n1377 ;
  assign n1380 = n1379 ^ n1374 ;
  assign n1385 = n1382 ^ n1380 ;
  assign n1368 = n1367 ^ n1365 ;
  assign n1386 = n1385 ^ n1368 ;
  assign n1340 = n1336 ^ n1334 ;
  assign n1341 = n1337 ^ n1335 ;
  assign n1342 = n1340 & n1341 ;
  assign n1344 = n1343 ^ n1342 ;
  assign n1345 = n1344 ^ n1339 ;
  assign n1350 = n1347 ^ n1345 ;
  assign n1333 = n1332 ^ n1330 ;
  assign n1351 = n1350 ^ n1333 ;
  assign n1436 = n1386 ^ n1351 ;
  assign n1459 = n1448 ^ n1436 ;
  assign n1460 = n1459 ^ n1293 ;
  assign n1507 = n1480 ^ n1460 ;
  assign n1001 = n990 ^ n970 ;
  assign n1508 = n1507 ^ n1001 ;
  assign n4415 = n2896 ^ n1508 ;
  assign n2784 = n2703 ^ n2695 ;
  assign n2785 = n2704 ^ n2696 ;
  assign n2795 = n2784 & n2785 ;
  assign n2782 = n2701 ^ n2693 ;
  assign n2783 = n2702 ^ n2694 ;
  assign n2794 = n2782 & n2783 ;
  assign n2799 = n2795 ^ n2794 ;
  assign n2780 = n2699 ^ n2691 ;
  assign n2781 = n2700 ^ n2692 ;
  assign n2787 = n2780 & n2781 ;
  assign n2778 = n2697 ^ n2689 ;
  assign n2779 = n2698 ^ n2690 ;
  assign n2786 = n2778 & n2779 ;
  assign n2791 = n2787 ^ n2786 ;
  assign n2815 = n2799 ^ n2791 ;
  assign n2825 = n2821 ^ n2815 ;
  assign n2826 = n2825 ^ n2772 ;
  assign n2849 = n2837 ^ n2826 ;
  assign n2685 = n2679 ^ n2670 ;
  assign n2850 = n2849 ^ n2685 ;
  assign n2897 = n2869 ^ n2850 ;
  assign n2382 = n2376 ^ n2364 ;
  assign n2390 = n2382 ^ n2359 ;
  assign n2898 = n2897 ^ n2390 ;
  assign n1396 = n1315 ^ n1307 ;
  assign n1397 = n1316 ^ n1308 ;
  assign n1407 = n1396 & n1397 ;
  assign n1394 = n1313 ^ n1305 ;
  assign n1395 = n1314 ^ n1306 ;
  assign n1406 = n1394 & n1395 ;
  assign n1411 = n1407 ^ n1406 ;
  assign n1392 = n1311 ^ n1303 ;
  assign n1393 = n1312 ^ n1304 ;
  assign n1399 = n1392 & n1393 ;
  assign n1390 = n1309 ^ n1301 ;
  assign n1391 = n1310 ^ n1302 ;
  assign n1398 = n1390 & n1391 ;
  assign n1403 = n1399 ^ n1398 ;
  assign n1427 = n1411 ^ n1403 ;
  assign n1437 = n1433 ^ n1427 ;
  assign n1438 = n1437 ^ n1384 ;
  assign n1461 = n1449 ^ n1438 ;
  assign n1297 = n1291 ^ n1282 ;
  assign n1462 = n1461 ^ n1297 ;
  assign n1509 = n1481 ^ n1462 ;
  assign n994 = n988 ^ n976 ;
  assign n1002 = n994 ^ n971 ;
  assign n1510 = n1509 ^ n1002 ;
  assign n4416 = n2898 ^ n1510 ;
  assign n2796 = n2784 ^ n2782 ;
  assign n2797 = n2785 ^ n2783 ;
  assign n2798 = n2796 & n2797 ;
  assign n2800 = n2799 ^ n2798 ;
  assign n2801 = n2800 ^ n2795 ;
  assign n2788 = n2780 ^ n2778 ;
  assign n2789 = n2781 ^ n2779 ;
  assign n2790 = n2788 & n2789 ;
  assign n2792 = n2791 ^ n2790 ;
  assign n2793 = n2792 ^ n2787 ;
  assign n2816 = n2801 ^ n2793 ;
  assign n2827 = n2822 ^ n2816 ;
  assign n2828 = n2827 ^ n2774 ;
  assign n2851 = n2838 ^ n2828 ;
  assign n2686 = n2681 ^ n2671 ;
  assign n2852 = n2851 ^ n2686 ;
  assign n2899 = n2870 ^ n2852 ;
  assign n2383 = n2378 ^ n2366 ;
  assign n2391 = n2383 ^ n2360 ;
  assign n2900 = n2899 ^ n2391 ;
  assign n1408 = n1396 ^ n1394 ;
  assign n1409 = n1397 ^ n1395 ;
  assign n1410 = n1408 & n1409 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1413 = n1412 ^ n1407 ;
  assign n1400 = n1392 ^ n1390 ;
  assign n1401 = n1393 ^ n1391 ;
  assign n1402 = n1400 & n1401 ;
  assign n1404 = n1403 ^ n1402 ;
  assign n1405 = n1404 ^ n1399 ;
  assign n1428 = n1413 ^ n1405 ;
  assign n1439 = n1434 ^ n1428 ;
  assign n1440 = n1439 ^ n1386 ;
  assign n1463 = n1450 ^ n1440 ;
  assign n1298 = n1293 ^ n1283 ;
  assign n1464 = n1463 ^ n1298 ;
  assign n1511 = n1482 ^ n1464 ;
  assign n995 = n990 ^ n978 ;
  assign n1003 = n995 ^ n972 ;
  assign n1512 = n1511 ^ n1003 ;
  assign n4417 = n2900 ^ n1512 ;
  assign n2805 = n2784 ^ n2780 ;
  assign n2806 = n2785 ^ n2781 ;
  assign n2808 = n2805 & n2806 ;
  assign n2803 = n2782 ^ n2778 ;
  assign n2804 = n2783 ^ n2779 ;
  assign n2807 = n2803 & n2804 ;
  assign n2812 = n2808 ^ n2807 ;
  assign n2817 = n2815 ^ n2812 ;
  assign n2818 = n2817 ^ n2801 ;
  assign n2829 = n2823 ^ n2818 ;
  assign n2776 = n2774 ^ n2769 ;
  assign n2830 = n2829 ^ n2776 ;
  assign n2853 = n2839 ^ n2830 ;
  assign n2683 = n2681 ^ n2675 ;
  assign n2687 = n2683 ^ n2672 ;
  assign n2854 = n2853 ^ n2687 ;
  assign n2901 = n2871 ^ n2854 ;
  assign n2380 = n2378 ^ n2372 ;
  assign n2384 = n2380 ^ n2368 ;
  assign n2392 = n2384 ^ n2361 ;
  assign n2902 = n2901 ^ n2392 ;
  assign n1417 = n1396 ^ n1392 ;
  assign n1418 = n1397 ^ n1393 ;
  assign n1420 = n1417 & n1418 ;
  assign n1415 = n1394 ^ n1390 ;
  assign n1416 = n1395 ^ n1391 ;
  assign n1419 = n1415 & n1416 ;
  assign n1424 = n1420 ^ n1419 ;
  assign n1429 = n1427 ^ n1424 ;
  assign n1430 = n1429 ^ n1413 ;
  assign n1441 = n1435 ^ n1430 ;
  assign n1388 = n1386 ^ n1381 ;
  assign n1442 = n1441 ^ n1388 ;
  assign n1465 = n1451 ^ n1442 ;
  assign n1295 = n1293 ^ n1287 ;
  assign n1299 = n1295 ^ n1284 ;
  assign n1466 = n1465 ^ n1299 ;
  assign n1513 = n1483 ^ n1466 ;
  assign n992 = n990 ^ n984 ;
  assign n996 = n992 ^ n980 ;
  assign n1004 = n996 ^ n973 ;
  assign n1514 = n1513 ^ n1004 ;
  assign n4418 = n2902 ^ n1514 ;
  assign n2809 = n2805 ^ n2803 ;
  assign n2810 = n2806 ^ n2804 ;
  assign n2811 = n2809 & n2810 ;
  assign n2813 = n2812 ^ n2811 ;
  assign n2814 = n2813 ^ n2808 ;
  assign n2819 = n2816 ^ n2814 ;
  assign n2802 = n2801 ^ n2799 ;
  assign n2820 = n2819 ^ n2802 ;
  assign n2831 = n2824 ^ n2820 ;
  assign n2775 = n2774 ^ n2772 ;
  assign n2777 = n2775 ^ n2770 ;
  assign n2832 = n2831 ^ n2777 ;
  assign n2855 = n2840 ^ n2832 ;
  assign n2682 = n2681 ^ n2679 ;
  assign n2684 = n2682 ^ n2677 ;
  assign n2688 = n2684 ^ n2673 ;
  assign n2856 = n2855 ^ n2688 ;
  assign n2903 = n2872 ^ n2856 ;
  assign n2379 = n2378 ^ n2376 ;
  assign n2381 = n2379 ^ n2374 ;
  assign n2385 = n2381 ^ n2370 ;
  assign n2393 = n2385 ^ n2362 ;
  assign n2904 = n2903 ^ n2393 ;
  assign n1421 = n1417 ^ n1415 ;
  assign n1422 = n1418 ^ n1416 ;
  assign n1423 = n1421 & n1422 ;
  assign n1425 = n1424 ^ n1423 ;
  assign n1426 = n1425 ^ n1420 ;
  assign n1431 = n1428 ^ n1426 ;
  assign n1414 = n1413 ^ n1411 ;
  assign n1432 = n1431 ^ n1414 ;
  assign n1443 = n1436 ^ n1432 ;
  assign n1387 = n1386 ^ n1384 ;
  assign n1389 = n1387 ^ n1382 ;
  assign n1444 = n1443 ^ n1389 ;
  assign n1467 = n1452 ^ n1444 ;
  assign n1294 = n1293 ^ n1291 ;
  assign n1296 = n1294 ^ n1289 ;
  assign n1300 = n1296 ^ n1285 ;
  assign n1468 = n1467 ^ n1300 ;
  assign n1515 = n1484 ^ n1468 ;
  assign n991 = n990 ^ n988 ;
  assign n993 = n991 ^ n986 ;
  assign n997 = n993 ^ n982 ;
  assign n1005 = n997 ^ n974 ;
  assign n1516 = n1515 ^ n1005 ;
  assign n4419 = n2904 ^ n1516 ;
  assign n2998 = x63 ^ x31 ;
  assign n2999 = x127 ^ x95 ;
  assign n3603 = n2998 & n2999 ;
  assign n2996 = x62 ^ x30 ;
  assign n2997 = x126 ^ x94 ;
  assign n3602 = n2996 & n2997 ;
  assign n3607 = n3603 ^ n3602 ;
  assign n2994 = x61 ^ x29 ;
  assign n2995 = x125 ^ x93 ;
  assign n3595 = n2994 & n2995 ;
  assign n2992 = x60 ^ x28 ;
  assign n2993 = x124 ^ x92 ;
  assign n3594 = n2992 & n2993 ;
  assign n3599 = n3595 ^ n3594 ;
  assign n3623 = n3607 ^ n3599 ;
  assign n2990 = x59 ^ x27 ;
  assign n2991 = x123 ^ x91 ;
  assign n3568 = n2990 & n2991 ;
  assign n2988 = x58 ^ x26 ;
  assign n2989 = x122 ^ x90 ;
  assign n3567 = n2988 & n2989 ;
  assign n3572 = n3568 ^ n3567 ;
  assign n2986 = x57 ^ x25 ;
  assign n2987 = x121 ^ x89 ;
  assign n3560 = n2986 & n2987 ;
  assign n2984 = x56 ^ x24 ;
  assign n2985 = x120 ^ x88 ;
  assign n3559 = n2984 & n2985 ;
  assign n3564 = n3560 ^ n3559 ;
  assign n3588 = n3572 ^ n3564 ;
  assign n3675 = n3623 ^ n3588 ;
  assign n2982 = x55 ^ x23 ;
  assign n2983 = x119 ^ x87 ;
  assign n3475 = n2982 & n2983 ;
  assign n2980 = x54 ^ x22 ;
  assign n2981 = x118 ^ x86 ;
  assign n3474 = n2980 & n2981 ;
  assign n3479 = n3475 ^ n3474 ;
  assign n2978 = x53 ^ x21 ;
  assign n2979 = x117 ^ x85 ;
  assign n3467 = n2978 & n2979 ;
  assign n2976 = x52 ^ x20 ;
  assign n2977 = x116 ^ x84 ;
  assign n3466 = n2976 & n2977 ;
  assign n3471 = n3467 ^ n3466 ;
  assign n3495 = n3479 ^ n3471 ;
  assign n2974 = x51 ^ x19 ;
  assign n2975 = x115 ^ x83 ;
  assign n3440 = n2974 & n2975 ;
  assign n2972 = x50 ^ x18 ;
  assign n2973 = x114 ^ x82 ;
  assign n3439 = n2972 & n2973 ;
  assign n3444 = n3440 ^ n3439 ;
  assign n2970 = x49 ^ x17 ;
  assign n2971 = x113 ^ x81 ;
  assign n3432 = n2970 & n2971 ;
  assign n2968 = x48 ^ x16 ;
  assign n2969 = x112 ^ x80 ;
  assign n3431 = n2968 & n2969 ;
  assign n3436 = n3432 ^ n3431 ;
  assign n3460 = n3444 ^ n3436 ;
  assign n3547 = n3495 ^ n3460 ;
  assign n3838 = n3675 ^ n3547 ;
  assign n2966 = x47 ^ x15 ;
  assign n2967 = x111 ^ x79 ;
  assign n3172 = n2966 & n2967 ;
  assign n2964 = x46 ^ x14 ;
  assign n2965 = x110 ^ x78 ;
  assign n3171 = n2964 & n2965 ;
  assign n3176 = n3172 ^ n3171 ;
  assign n2962 = x45 ^ x13 ;
  assign n2963 = x109 ^ x77 ;
  assign n3164 = n2962 & n2963 ;
  assign n2960 = x44 ^ x12 ;
  assign n2961 = x108 ^ x76 ;
  assign n3163 = n2960 & n2961 ;
  assign n3168 = n3164 ^ n3163 ;
  assign n3192 = n3176 ^ n3168 ;
  assign n2958 = x43 ^ x11 ;
  assign n2959 = x107 ^ x75 ;
  assign n3137 = n2958 & n2959 ;
  assign n2956 = x42 ^ x10 ;
  assign n2957 = x106 ^ x74 ;
  assign n3136 = n2956 & n2957 ;
  assign n3141 = n3137 ^ n3136 ;
  assign n2954 = x41 ^ x9 ;
  assign n2955 = x105 ^ x73 ;
  assign n3129 = n2954 & n2955 ;
  assign n2952 = x40 ^ x8 ;
  assign n2953 = x104 ^ x72 ;
  assign n3128 = n2952 & n2953 ;
  assign n3133 = n3129 ^ n3128 ;
  assign n3157 = n3141 ^ n3133 ;
  assign n3244 = n3192 ^ n3157 ;
  assign n2950 = x39 ^ x7 ;
  assign n2951 = x103 ^ x71 ;
  assign n3044 = n2950 & n2951 ;
  assign n2948 = x38 ^ x6 ;
  assign n2949 = x102 ^ x70 ;
  assign n3043 = n2948 & n2949 ;
  assign n3048 = n3044 ^ n3043 ;
  assign n2946 = x37 ^ x5 ;
  assign n2947 = x101 ^ x69 ;
  assign n3036 = n2946 & n2947 ;
  assign n2944 = x36 ^ x4 ;
  assign n2945 = x100 ^ x68 ;
  assign n3035 = n2944 & n2945 ;
  assign n3040 = n3036 ^ n3035 ;
  assign n3064 = n3048 ^ n3040 ;
  assign n2942 = x35 ^ x3 ;
  assign n2943 = x99 ^ x67 ;
  assign n3009 = n2942 & n2943 ;
  assign n2940 = x34 ^ x2 ;
  assign n2941 = x98 ^ x66 ;
  assign n3008 = n2940 & n2941 ;
  assign n3013 = n3009 ^ n3008 ;
  assign n2938 = x33 ^ x1 ;
  assign n2939 = x97 ^ x65 ;
  assign n3001 = n2938 & n2939 ;
  assign n2936 = x32 ^ x0 ;
  assign n2937 = x96 ^ x64 ;
  assign n3000 = n2936 & n2937 ;
  assign n3005 = n3001 ^ n3000 ;
  assign n3029 = n3013 ^ n3005 ;
  assign n3116 = n3064 ^ n3029 ;
  assign n3407 = n3244 ^ n3116 ;
  assign n4340 = n3838 ^ n3407 ;
  assign n4420 = n4388 ^ n4340 ;
  assign n4421 = n4420 ^ n2874 ;
  assign n3604 = n2998 ^ n2996 ;
  assign n3605 = n2999 ^ n2997 ;
  assign n3606 = n3604 & n3605 ;
  assign n3608 = n3607 ^ n3606 ;
  assign n3609 = n3608 ^ n3603 ;
  assign n3596 = n2994 ^ n2992 ;
  assign n3597 = n2995 ^ n2993 ;
  assign n3598 = n3596 & n3597 ;
  assign n3600 = n3599 ^ n3598 ;
  assign n3601 = n3600 ^ n3595 ;
  assign n3624 = n3609 ^ n3601 ;
  assign n3569 = n2990 ^ n2988 ;
  assign n3570 = n2991 ^ n2989 ;
  assign n3571 = n3569 & n3570 ;
  assign n3573 = n3572 ^ n3571 ;
  assign n3574 = n3573 ^ n3568 ;
  assign n3561 = n2986 ^ n2984 ;
  assign n3562 = n2987 ^ n2985 ;
  assign n3563 = n3561 & n3562 ;
  assign n3565 = n3564 ^ n3563 ;
  assign n3566 = n3565 ^ n3560 ;
  assign n3589 = n3574 ^ n3566 ;
  assign n3676 = n3624 ^ n3589 ;
  assign n3476 = n2982 ^ n2980 ;
  assign n3477 = n2983 ^ n2981 ;
  assign n3478 = n3476 & n3477 ;
  assign n3480 = n3479 ^ n3478 ;
  assign n3481 = n3480 ^ n3475 ;
  assign n3468 = n2978 ^ n2976 ;
  assign n3469 = n2979 ^ n2977 ;
  assign n3470 = n3468 & n3469 ;
  assign n3472 = n3471 ^ n3470 ;
  assign n3473 = n3472 ^ n3467 ;
  assign n3496 = n3481 ^ n3473 ;
  assign n3441 = n2974 ^ n2972 ;
  assign n3442 = n2975 ^ n2973 ;
  assign n3443 = n3441 & n3442 ;
  assign n3445 = n3444 ^ n3443 ;
  assign n3446 = n3445 ^ n3440 ;
  assign n3433 = n2970 ^ n2968 ;
  assign n3434 = n2971 ^ n2969 ;
  assign n3435 = n3433 & n3434 ;
  assign n3437 = n3436 ^ n3435 ;
  assign n3438 = n3437 ^ n3432 ;
  assign n3461 = n3446 ^ n3438 ;
  assign n3548 = n3496 ^ n3461 ;
  assign n3839 = n3676 ^ n3548 ;
  assign n3173 = n2966 ^ n2964 ;
  assign n3174 = n2967 ^ n2965 ;
  assign n3175 = n3173 & n3174 ;
  assign n3177 = n3176 ^ n3175 ;
  assign n3178 = n3177 ^ n3172 ;
  assign n3165 = n2962 ^ n2960 ;
  assign n3166 = n2963 ^ n2961 ;
  assign n3167 = n3165 & n3166 ;
  assign n3169 = n3168 ^ n3167 ;
  assign n3170 = n3169 ^ n3164 ;
  assign n3193 = n3178 ^ n3170 ;
  assign n3138 = n2958 ^ n2956 ;
  assign n3139 = n2959 ^ n2957 ;
  assign n3140 = n3138 & n3139 ;
  assign n3142 = n3141 ^ n3140 ;
  assign n3143 = n3142 ^ n3137 ;
  assign n3130 = n2954 ^ n2952 ;
  assign n3131 = n2955 ^ n2953 ;
  assign n3132 = n3130 & n3131 ;
  assign n3134 = n3133 ^ n3132 ;
  assign n3135 = n3134 ^ n3129 ;
  assign n3158 = n3143 ^ n3135 ;
  assign n3245 = n3193 ^ n3158 ;
  assign n3045 = n2950 ^ n2948 ;
  assign n3046 = n2951 ^ n2949 ;
  assign n3047 = n3045 & n3046 ;
  assign n3049 = n3048 ^ n3047 ;
  assign n3050 = n3049 ^ n3044 ;
  assign n3037 = n2946 ^ n2944 ;
  assign n3038 = n2947 ^ n2945 ;
  assign n3039 = n3037 & n3038 ;
  assign n3041 = n3040 ^ n3039 ;
  assign n3042 = n3041 ^ n3036 ;
  assign n3065 = n3050 ^ n3042 ;
  assign n3010 = n2942 ^ n2940 ;
  assign n3011 = n2943 ^ n2941 ;
  assign n3012 = n3010 & n3011 ;
  assign n3014 = n3013 ^ n3012 ;
  assign n3015 = n3014 ^ n3009 ;
  assign n3002 = n2938 ^ n2936 ;
  assign n3003 = n2939 ^ n2937 ;
  assign n3004 = n3002 & n3003 ;
  assign n3006 = n3005 ^ n3004 ;
  assign n3007 = n3006 ^ n3001 ;
  assign n3030 = n3015 ^ n3007 ;
  assign n3117 = n3065 ^ n3030 ;
  assign n3408 = n3245 ^ n3117 ;
  assign n4341 = n3839 ^ n3408 ;
  assign n4422 = n4389 ^ n4341 ;
  assign n4423 = n4422 ^ n2876 ;
  assign n3613 = n2998 ^ n2994 ;
  assign n3614 = n2999 ^ n2995 ;
  assign n3616 = n3613 & n3614 ;
  assign n3611 = n2996 ^ n2992 ;
  assign n3612 = n2997 ^ n2993 ;
  assign n3615 = n3611 & n3612 ;
  assign n3620 = n3616 ^ n3615 ;
  assign n3625 = n3623 ^ n3620 ;
  assign n3626 = n3625 ^ n3609 ;
  assign n3578 = n2990 ^ n2986 ;
  assign n3579 = n2991 ^ n2987 ;
  assign n3581 = n3578 & n3579 ;
  assign n3576 = n2988 ^ n2984 ;
  assign n3577 = n2989 ^ n2985 ;
  assign n3580 = n3576 & n3577 ;
  assign n3585 = n3581 ^ n3580 ;
  assign n3590 = n3588 ^ n3585 ;
  assign n3591 = n3590 ^ n3574 ;
  assign n3677 = n3626 ^ n3591 ;
  assign n3485 = n2982 ^ n2978 ;
  assign n3486 = n2983 ^ n2979 ;
  assign n3488 = n3485 & n3486 ;
  assign n3483 = n2980 ^ n2976 ;
  assign n3484 = n2981 ^ n2977 ;
  assign n3487 = n3483 & n3484 ;
  assign n3492 = n3488 ^ n3487 ;
  assign n3497 = n3495 ^ n3492 ;
  assign n3498 = n3497 ^ n3481 ;
  assign n3450 = n2974 ^ n2970 ;
  assign n3451 = n2975 ^ n2971 ;
  assign n3453 = n3450 & n3451 ;
  assign n3448 = n2972 ^ n2968 ;
  assign n3449 = n2973 ^ n2969 ;
  assign n3452 = n3448 & n3449 ;
  assign n3457 = n3453 ^ n3452 ;
  assign n3462 = n3460 ^ n3457 ;
  assign n3463 = n3462 ^ n3446 ;
  assign n3549 = n3498 ^ n3463 ;
  assign n3840 = n3677 ^ n3549 ;
  assign n3182 = n2966 ^ n2962 ;
  assign n3183 = n2967 ^ n2963 ;
  assign n3185 = n3182 & n3183 ;
  assign n3180 = n2964 ^ n2960 ;
  assign n3181 = n2965 ^ n2961 ;
  assign n3184 = n3180 & n3181 ;
  assign n3189 = n3185 ^ n3184 ;
  assign n3194 = n3192 ^ n3189 ;
  assign n3195 = n3194 ^ n3178 ;
  assign n3147 = n2958 ^ n2954 ;
  assign n3148 = n2959 ^ n2955 ;
  assign n3150 = n3147 & n3148 ;
  assign n3145 = n2956 ^ n2952 ;
  assign n3146 = n2957 ^ n2953 ;
  assign n3149 = n3145 & n3146 ;
  assign n3154 = n3150 ^ n3149 ;
  assign n3159 = n3157 ^ n3154 ;
  assign n3160 = n3159 ^ n3143 ;
  assign n3246 = n3195 ^ n3160 ;
  assign n3054 = n2950 ^ n2946 ;
  assign n3055 = n2951 ^ n2947 ;
  assign n3057 = n3054 & n3055 ;
  assign n3052 = n2948 ^ n2944 ;
  assign n3053 = n2949 ^ n2945 ;
  assign n3056 = n3052 & n3053 ;
  assign n3061 = n3057 ^ n3056 ;
  assign n3066 = n3064 ^ n3061 ;
  assign n3067 = n3066 ^ n3050 ;
  assign n3019 = n2942 ^ n2938 ;
  assign n3020 = n2943 ^ n2939 ;
  assign n3022 = n3019 & n3020 ;
  assign n3017 = n2940 ^ n2936 ;
  assign n3018 = n2941 ^ n2937 ;
  assign n3021 = n3017 & n3018 ;
  assign n3026 = n3022 ^ n3021 ;
  assign n3031 = n3029 ^ n3026 ;
  assign n3032 = n3031 ^ n3015 ;
  assign n3118 = n3067 ^ n3032 ;
  assign n3409 = n3246 ^ n3118 ;
  assign n4342 = n3840 ^ n3409 ;
  assign n4424 = n4390 ^ n4342 ;
  assign n4425 = n4424 ^ n2878 ;
  assign n3617 = n3613 ^ n3611 ;
  assign n3618 = n3614 ^ n3612 ;
  assign n3619 = n3617 & n3618 ;
  assign n3621 = n3620 ^ n3619 ;
  assign n3622 = n3621 ^ n3616 ;
  assign n3627 = n3624 ^ n3622 ;
  assign n3610 = n3609 ^ n3607 ;
  assign n3628 = n3627 ^ n3610 ;
  assign n3582 = n3578 ^ n3576 ;
  assign n3583 = n3579 ^ n3577 ;
  assign n3584 = n3582 & n3583 ;
  assign n3586 = n3585 ^ n3584 ;
  assign n3587 = n3586 ^ n3581 ;
  assign n3592 = n3589 ^ n3587 ;
  assign n3575 = n3574 ^ n3572 ;
  assign n3593 = n3592 ^ n3575 ;
  assign n3678 = n3628 ^ n3593 ;
  assign n3489 = n3485 ^ n3483 ;
  assign n3490 = n3486 ^ n3484 ;
  assign n3491 = n3489 & n3490 ;
  assign n3493 = n3492 ^ n3491 ;
  assign n3494 = n3493 ^ n3488 ;
  assign n3499 = n3496 ^ n3494 ;
  assign n3482 = n3481 ^ n3479 ;
  assign n3500 = n3499 ^ n3482 ;
  assign n3454 = n3450 ^ n3448 ;
  assign n3455 = n3451 ^ n3449 ;
  assign n3456 = n3454 & n3455 ;
  assign n3458 = n3457 ^ n3456 ;
  assign n3459 = n3458 ^ n3453 ;
  assign n3464 = n3461 ^ n3459 ;
  assign n3447 = n3446 ^ n3444 ;
  assign n3465 = n3464 ^ n3447 ;
  assign n3550 = n3500 ^ n3465 ;
  assign n3841 = n3678 ^ n3550 ;
  assign n3186 = n3182 ^ n3180 ;
  assign n3187 = n3183 ^ n3181 ;
  assign n3188 = n3186 & n3187 ;
  assign n3190 = n3189 ^ n3188 ;
  assign n3191 = n3190 ^ n3185 ;
  assign n3196 = n3193 ^ n3191 ;
  assign n3179 = n3178 ^ n3176 ;
  assign n3197 = n3196 ^ n3179 ;
  assign n3151 = n3147 ^ n3145 ;
  assign n3152 = n3148 ^ n3146 ;
  assign n3153 = n3151 & n3152 ;
  assign n3155 = n3154 ^ n3153 ;
  assign n3156 = n3155 ^ n3150 ;
  assign n3161 = n3158 ^ n3156 ;
  assign n3144 = n3143 ^ n3141 ;
  assign n3162 = n3161 ^ n3144 ;
  assign n3247 = n3197 ^ n3162 ;
  assign n3058 = n3054 ^ n3052 ;
  assign n3059 = n3055 ^ n3053 ;
  assign n3060 = n3058 & n3059 ;
  assign n3062 = n3061 ^ n3060 ;
  assign n3063 = n3062 ^ n3057 ;
  assign n3068 = n3065 ^ n3063 ;
  assign n3051 = n3050 ^ n3048 ;
  assign n3069 = n3068 ^ n3051 ;
  assign n3023 = n3019 ^ n3017 ;
  assign n3024 = n3020 ^ n3018 ;
  assign n3025 = n3023 & n3024 ;
  assign n3027 = n3026 ^ n3025 ;
  assign n3028 = n3027 ^ n3022 ;
  assign n3033 = n3030 ^ n3028 ;
  assign n3016 = n3015 ^ n3013 ;
  assign n3034 = n3033 ^ n3016 ;
  assign n3119 = n3069 ^ n3034 ;
  assign n3410 = n3247 ^ n3119 ;
  assign n4343 = n3841 ^ n3410 ;
  assign n4426 = n4391 ^ n4343 ;
  assign n4427 = n4426 ^ n2880 ;
  assign n3638 = n2998 ^ n2990 ;
  assign n3639 = n2999 ^ n2991 ;
  assign n3649 = n3638 & n3639 ;
  assign n3636 = n2996 ^ n2988 ;
  assign n3637 = n2997 ^ n2989 ;
  assign n3648 = n3636 & n3637 ;
  assign n3653 = n3649 ^ n3648 ;
  assign n3634 = n2994 ^ n2986 ;
  assign n3635 = n2995 ^ n2987 ;
  assign n3641 = n3634 & n3635 ;
  assign n3632 = n2992 ^ n2984 ;
  assign n3633 = n2993 ^ n2985 ;
  assign n3640 = n3632 & n3633 ;
  assign n3645 = n3641 ^ n3640 ;
  assign n3669 = n3653 ^ n3645 ;
  assign n3679 = n3675 ^ n3669 ;
  assign n3680 = n3679 ^ n3626 ;
  assign n3510 = n2982 ^ n2974 ;
  assign n3511 = n2983 ^ n2975 ;
  assign n3521 = n3510 & n3511 ;
  assign n3508 = n2980 ^ n2972 ;
  assign n3509 = n2981 ^ n2973 ;
  assign n3520 = n3508 & n3509 ;
  assign n3525 = n3521 ^ n3520 ;
  assign n3506 = n2978 ^ n2970 ;
  assign n3507 = n2979 ^ n2971 ;
  assign n3513 = n3506 & n3507 ;
  assign n3504 = n2976 ^ n2968 ;
  assign n3505 = n2977 ^ n2969 ;
  assign n3512 = n3504 & n3505 ;
  assign n3517 = n3513 ^ n3512 ;
  assign n3541 = n3525 ^ n3517 ;
  assign n3551 = n3547 ^ n3541 ;
  assign n3552 = n3551 ^ n3498 ;
  assign n3842 = n3680 ^ n3552 ;
  assign n3207 = n2966 ^ n2958 ;
  assign n3208 = n2967 ^ n2959 ;
  assign n3218 = n3207 & n3208 ;
  assign n3205 = n2964 ^ n2956 ;
  assign n3206 = n2965 ^ n2957 ;
  assign n3217 = n3205 & n3206 ;
  assign n3222 = n3218 ^ n3217 ;
  assign n3203 = n2962 ^ n2954 ;
  assign n3204 = n2963 ^ n2955 ;
  assign n3210 = n3203 & n3204 ;
  assign n3201 = n2960 ^ n2952 ;
  assign n3202 = n2961 ^ n2953 ;
  assign n3209 = n3201 & n3202 ;
  assign n3214 = n3210 ^ n3209 ;
  assign n3238 = n3222 ^ n3214 ;
  assign n3248 = n3244 ^ n3238 ;
  assign n3249 = n3248 ^ n3195 ;
  assign n3079 = n2950 ^ n2942 ;
  assign n3080 = n2951 ^ n2943 ;
  assign n3090 = n3079 & n3080 ;
  assign n3077 = n2948 ^ n2940 ;
  assign n3078 = n2949 ^ n2941 ;
  assign n3089 = n3077 & n3078 ;
  assign n3094 = n3090 ^ n3089 ;
  assign n3075 = n2946 ^ n2938 ;
  assign n3076 = n2947 ^ n2939 ;
  assign n3082 = n3075 & n3076 ;
  assign n3073 = n2944 ^ n2936 ;
  assign n3074 = n2945 ^ n2937 ;
  assign n3081 = n3073 & n3074 ;
  assign n3086 = n3082 ^ n3081 ;
  assign n3110 = n3094 ^ n3086 ;
  assign n3120 = n3116 ^ n3110 ;
  assign n3121 = n3120 ^ n3067 ;
  assign n3411 = n3249 ^ n3121 ;
  assign n4344 = n3842 ^ n3411 ;
  assign n4428 = n4392 ^ n4344 ;
  assign n4429 = n4428 ^ n2882 ;
  assign n3650 = n3638 ^ n3636 ;
  assign n3651 = n3639 ^ n3637 ;
  assign n3652 = n3650 & n3651 ;
  assign n3654 = n3653 ^ n3652 ;
  assign n3655 = n3654 ^ n3649 ;
  assign n3642 = n3634 ^ n3632 ;
  assign n3643 = n3635 ^ n3633 ;
  assign n3644 = n3642 & n3643 ;
  assign n3646 = n3645 ^ n3644 ;
  assign n3647 = n3646 ^ n3641 ;
  assign n3670 = n3655 ^ n3647 ;
  assign n3681 = n3676 ^ n3670 ;
  assign n3682 = n3681 ^ n3628 ;
  assign n3522 = n3510 ^ n3508 ;
  assign n3523 = n3511 ^ n3509 ;
  assign n3524 = n3522 & n3523 ;
  assign n3526 = n3525 ^ n3524 ;
  assign n3527 = n3526 ^ n3521 ;
  assign n3514 = n3506 ^ n3504 ;
  assign n3515 = n3507 ^ n3505 ;
  assign n3516 = n3514 & n3515 ;
  assign n3518 = n3517 ^ n3516 ;
  assign n3519 = n3518 ^ n3513 ;
  assign n3542 = n3527 ^ n3519 ;
  assign n3553 = n3548 ^ n3542 ;
  assign n3554 = n3553 ^ n3500 ;
  assign n3843 = n3682 ^ n3554 ;
  assign n3219 = n3207 ^ n3205 ;
  assign n3220 = n3208 ^ n3206 ;
  assign n3221 = n3219 & n3220 ;
  assign n3223 = n3222 ^ n3221 ;
  assign n3224 = n3223 ^ n3218 ;
  assign n3211 = n3203 ^ n3201 ;
  assign n3212 = n3204 ^ n3202 ;
  assign n3213 = n3211 & n3212 ;
  assign n3215 = n3214 ^ n3213 ;
  assign n3216 = n3215 ^ n3210 ;
  assign n3239 = n3224 ^ n3216 ;
  assign n3250 = n3245 ^ n3239 ;
  assign n3251 = n3250 ^ n3197 ;
  assign n3091 = n3079 ^ n3077 ;
  assign n3092 = n3080 ^ n3078 ;
  assign n3093 = n3091 & n3092 ;
  assign n3095 = n3094 ^ n3093 ;
  assign n3096 = n3095 ^ n3090 ;
  assign n3083 = n3075 ^ n3073 ;
  assign n3084 = n3076 ^ n3074 ;
  assign n3085 = n3083 & n3084 ;
  assign n3087 = n3086 ^ n3085 ;
  assign n3088 = n3087 ^ n3082 ;
  assign n3111 = n3096 ^ n3088 ;
  assign n3122 = n3117 ^ n3111 ;
  assign n3123 = n3122 ^ n3069 ;
  assign n3412 = n3251 ^ n3123 ;
  assign n4345 = n3843 ^ n3412 ;
  assign n4430 = n4393 ^ n4345 ;
  assign n4431 = n4430 ^ n2884 ;
  assign n3659 = n3638 ^ n3634 ;
  assign n3660 = n3639 ^ n3635 ;
  assign n3662 = n3659 & n3660 ;
  assign n3657 = n3636 ^ n3632 ;
  assign n3658 = n3637 ^ n3633 ;
  assign n3661 = n3657 & n3658 ;
  assign n3666 = n3662 ^ n3661 ;
  assign n3671 = n3669 ^ n3666 ;
  assign n3672 = n3671 ^ n3655 ;
  assign n3683 = n3677 ^ n3672 ;
  assign n3630 = n3628 ^ n3623 ;
  assign n3684 = n3683 ^ n3630 ;
  assign n3531 = n3510 ^ n3506 ;
  assign n3532 = n3511 ^ n3507 ;
  assign n3534 = n3531 & n3532 ;
  assign n3529 = n3508 ^ n3504 ;
  assign n3530 = n3509 ^ n3505 ;
  assign n3533 = n3529 & n3530 ;
  assign n3538 = n3534 ^ n3533 ;
  assign n3543 = n3541 ^ n3538 ;
  assign n3544 = n3543 ^ n3527 ;
  assign n3555 = n3549 ^ n3544 ;
  assign n3502 = n3500 ^ n3495 ;
  assign n3556 = n3555 ^ n3502 ;
  assign n3844 = n3684 ^ n3556 ;
  assign n3228 = n3207 ^ n3203 ;
  assign n3229 = n3208 ^ n3204 ;
  assign n3231 = n3228 & n3229 ;
  assign n3226 = n3205 ^ n3201 ;
  assign n3227 = n3206 ^ n3202 ;
  assign n3230 = n3226 & n3227 ;
  assign n3235 = n3231 ^ n3230 ;
  assign n3240 = n3238 ^ n3235 ;
  assign n3241 = n3240 ^ n3224 ;
  assign n3252 = n3246 ^ n3241 ;
  assign n3199 = n3197 ^ n3192 ;
  assign n3253 = n3252 ^ n3199 ;
  assign n3100 = n3079 ^ n3075 ;
  assign n3101 = n3080 ^ n3076 ;
  assign n3103 = n3100 & n3101 ;
  assign n3098 = n3077 ^ n3073 ;
  assign n3099 = n3078 ^ n3074 ;
  assign n3102 = n3098 & n3099 ;
  assign n3107 = n3103 ^ n3102 ;
  assign n3112 = n3110 ^ n3107 ;
  assign n3113 = n3112 ^ n3096 ;
  assign n3124 = n3118 ^ n3113 ;
  assign n3071 = n3069 ^ n3064 ;
  assign n3125 = n3124 ^ n3071 ;
  assign n3413 = n3253 ^ n3125 ;
  assign n4346 = n3844 ^ n3413 ;
  assign n4432 = n4394 ^ n4346 ;
  assign n4433 = n4432 ^ n2886 ;
  assign n3663 = n3659 ^ n3657 ;
  assign n3664 = n3660 ^ n3658 ;
  assign n3665 = n3663 & n3664 ;
  assign n3667 = n3666 ^ n3665 ;
  assign n3668 = n3667 ^ n3662 ;
  assign n3673 = n3670 ^ n3668 ;
  assign n3656 = n3655 ^ n3653 ;
  assign n3674 = n3673 ^ n3656 ;
  assign n3685 = n3678 ^ n3674 ;
  assign n3629 = n3628 ^ n3626 ;
  assign n3631 = n3629 ^ n3624 ;
  assign n3686 = n3685 ^ n3631 ;
  assign n3535 = n3531 ^ n3529 ;
  assign n3536 = n3532 ^ n3530 ;
  assign n3537 = n3535 & n3536 ;
  assign n3539 = n3538 ^ n3537 ;
  assign n3540 = n3539 ^ n3534 ;
  assign n3545 = n3542 ^ n3540 ;
  assign n3528 = n3527 ^ n3525 ;
  assign n3546 = n3545 ^ n3528 ;
  assign n3557 = n3550 ^ n3546 ;
  assign n3501 = n3500 ^ n3498 ;
  assign n3503 = n3501 ^ n3496 ;
  assign n3558 = n3557 ^ n3503 ;
  assign n3845 = n3686 ^ n3558 ;
  assign n3232 = n3228 ^ n3226 ;
  assign n3233 = n3229 ^ n3227 ;
  assign n3234 = n3232 & n3233 ;
  assign n3236 = n3235 ^ n3234 ;
  assign n3237 = n3236 ^ n3231 ;
  assign n3242 = n3239 ^ n3237 ;
  assign n3225 = n3224 ^ n3222 ;
  assign n3243 = n3242 ^ n3225 ;
  assign n3254 = n3247 ^ n3243 ;
  assign n3198 = n3197 ^ n3195 ;
  assign n3200 = n3198 ^ n3193 ;
  assign n3255 = n3254 ^ n3200 ;
  assign n3104 = n3100 ^ n3098 ;
  assign n3105 = n3101 ^ n3099 ;
  assign n3106 = n3104 & n3105 ;
  assign n3108 = n3107 ^ n3106 ;
  assign n3109 = n3108 ^ n3103 ;
  assign n3114 = n3111 ^ n3109 ;
  assign n3097 = n3096 ^ n3094 ;
  assign n3115 = n3114 ^ n3097 ;
  assign n3126 = n3119 ^ n3115 ;
  assign n3070 = n3069 ^ n3067 ;
  assign n3072 = n3070 ^ n3065 ;
  assign n3127 = n3126 ^ n3072 ;
  assign n3414 = n3255 ^ n3127 ;
  assign n4347 = n3845 ^ n3414 ;
  assign n4434 = n4395 ^ n4347 ;
  assign n4435 = n4434 ^ n2888 ;
  assign n3708 = n2998 ^ n2982 ;
  assign n3709 = n2999 ^ n2983 ;
  assign n3754 = n3708 & n3709 ;
  assign n3706 = n2996 ^ n2980 ;
  assign n3707 = n2997 ^ n2981 ;
  assign n3753 = n3706 & n3707 ;
  assign n3758 = n3754 ^ n3753 ;
  assign n3704 = n2994 ^ n2978 ;
  assign n3705 = n2995 ^ n2979 ;
  assign n3746 = n3704 & n3705 ;
  assign n3702 = n2992 ^ n2976 ;
  assign n3703 = n2993 ^ n2977 ;
  assign n3745 = n3702 & n3703 ;
  assign n3750 = n3746 ^ n3745 ;
  assign n3774 = n3758 ^ n3750 ;
  assign n3700 = n2990 ^ n2974 ;
  assign n3701 = n2991 ^ n2975 ;
  assign n3719 = n3700 & n3701 ;
  assign n3698 = n2988 ^ n2972 ;
  assign n3699 = n2989 ^ n2973 ;
  assign n3718 = n3698 & n3699 ;
  assign n3723 = n3719 ^ n3718 ;
  assign n3696 = n2986 ^ n2970 ;
  assign n3697 = n2987 ^ n2971 ;
  assign n3711 = n3696 & n3697 ;
  assign n3694 = n2984 ^ n2968 ;
  assign n3695 = n2985 ^ n2969 ;
  assign n3710 = n3694 & n3695 ;
  assign n3715 = n3711 ^ n3710 ;
  assign n3739 = n3723 ^ n3715 ;
  assign n3826 = n3774 ^ n3739 ;
  assign n3846 = n3838 ^ n3826 ;
  assign n3847 = n3846 ^ n3680 ;
  assign n3277 = n2966 ^ n2950 ;
  assign n3278 = n2967 ^ n2951 ;
  assign n3323 = n3277 & n3278 ;
  assign n3275 = n2964 ^ n2948 ;
  assign n3276 = n2965 ^ n2949 ;
  assign n3322 = n3275 & n3276 ;
  assign n3327 = n3323 ^ n3322 ;
  assign n3273 = n2962 ^ n2946 ;
  assign n3274 = n2963 ^ n2947 ;
  assign n3315 = n3273 & n3274 ;
  assign n3271 = n2960 ^ n2944 ;
  assign n3272 = n2961 ^ n2945 ;
  assign n3314 = n3271 & n3272 ;
  assign n3319 = n3315 ^ n3314 ;
  assign n3343 = n3327 ^ n3319 ;
  assign n3269 = n2958 ^ n2942 ;
  assign n3270 = n2959 ^ n2943 ;
  assign n3288 = n3269 & n3270 ;
  assign n3267 = n2956 ^ n2940 ;
  assign n3268 = n2957 ^ n2941 ;
  assign n3287 = n3267 & n3268 ;
  assign n3292 = n3288 ^ n3287 ;
  assign n3265 = n2954 ^ n2938 ;
  assign n3266 = n2955 ^ n2939 ;
  assign n3280 = n3265 & n3266 ;
  assign n3263 = n2952 ^ n2936 ;
  assign n3264 = n2953 ^ n2937 ;
  assign n3279 = n3263 & n3264 ;
  assign n3284 = n3280 ^ n3279 ;
  assign n3308 = n3292 ^ n3284 ;
  assign n3395 = n3343 ^ n3308 ;
  assign n3415 = n3407 ^ n3395 ;
  assign n3416 = n3415 ^ n3249 ;
  assign n4348 = n3847 ^ n3416 ;
  assign n4436 = n4396 ^ n4348 ;
  assign n4437 = n4436 ^ n2890 ;
  assign n3755 = n3708 ^ n3706 ;
  assign n3756 = n3709 ^ n3707 ;
  assign n3757 = n3755 & n3756 ;
  assign n3759 = n3758 ^ n3757 ;
  assign n3760 = n3759 ^ n3754 ;
  assign n3747 = n3704 ^ n3702 ;
  assign n3748 = n3705 ^ n3703 ;
  assign n3749 = n3747 & n3748 ;
  assign n3751 = n3750 ^ n3749 ;
  assign n3752 = n3751 ^ n3746 ;
  assign n3775 = n3760 ^ n3752 ;
  assign n3720 = n3700 ^ n3698 ;
  assign n3721 = n3701 ^ n3699 ;
  assign n3722 = n3720 & n3721 ;
  assign n3724 = n3723 ^ n3722 ;
  assign n3725 = n3724 ^ n3719 ;
  assign n3712 = n3696 ^ n3694 ;
  assign n3713 = n3697 ^ n3695 ;
  assign n3714 = n3712 & n3713 ;
  assign n3716 = n3715 ^ n3714 ;
  assign n3717 = n3716 ^ n3711 ;
  assign n3740 = n3725 ^ n3717 ;
  assign n3827 = n3775 ^ n3740 ;
  assign n3848 = n3839 ^ n3827 ;
  assign n3849 = n3848 ^ n3682 ;
  assign n3324 = n3277 ^ n3275 ;
  assign n3325 = n3278 ^ n3276 ;
  assign n3326 = n3324 & n3325 ;
  assign n3328 = n3327 ^ n3326 ;
  assign n3329 = n3328 ^ n3323 ;
  assign n3316 = n3273 ^ n3271 ;
  assign n3317 = n3274 ^ n3272 ;
  assign n3318 = n3316 & n3317 ;
  assign n3320 = n3319 ^ n3318 ;
  assign n3321 = n3320 ^ n3315 ;
  assign n3344 = n3329 ^ n3321 ;
  assign n3289 = n3269 ^ n3267 ;
  assign n3290 = n3270 ^ n3268 ;
  assign n3291 = n3289 & n3290 ;
  assign n3293 = n3292 ^ n3291 ;
  assign n3294 = n3293 ^ n3288 ;
  assign n3281 = n3265 ^ n3263 ;
  assign n3282 = n3266 ^ n3264 ;
  assign n3283 = n3281 & n3282 ;
  assign n3285 = n3284 ^ n3283 ;
  assign n3286 = n3285 ^ n3280 ;
  assign n3309 = n3294 ^ n3286 ;
  assign n3396 = n3344 ^ n3309 ;
  assign n3417 = n3408 ^ n3396 ;
  assign n3418 = n3417 ^ n3251 ;
  assign n4349 = n3849 ^ n3418 ;
  assign n4438 = n4397 ^ n4349 ;
  assign n4439 = n4438 ^ n2892 ;
  assign n3764 = n3708 ^ n3704 ;
  assign n3765 = n3709 ^ n3705 ;
  assign n3767 = n3764 & n3765 ;
  assign n3762 = n3706 ^ n3702 ;
  assign n3763 = n3707 ^ n3703 ;
  assign n3766 = n3762 & n3763 ;
  assign n3771 = n3767 ^ n3766 ;
  assign n3776 = n3774 ^ n3771 ;
  assign n3777 = n3776 ^ n3760 ;
  assign n3729 = n3700 ^ n3696 ;
  assign n3730 = n3701 ^ n3697 ;
  assign n3732 = n3729 & n3730 ;
  assign n3727 = n3698 ^ n3694 ;
  assign n3728 = n3699 ^ n3695 ;
  assign n3731 = n3727 & n3728 ;
  assign n3736 = n3732 ^ n3731 ;
  assign n3741 = n3739 ^ n3736 ;
  assign n3742 = n3741 ^ n3725 ;
  assign n3828 = n3777 ^ n3742 ;
  assign n3850 = n3840 ^ n3828 ;
  assign n3851 = n3850 ^ n3684 ;
  assign n3333 = n3277 ^ n3273 ;
  assign n3334 = n3278 ^ n3274 ;
  assign n3336 = n3333 & n3334 ;
  assign n3331 = n3275 ^ n3271 ;
  assign n3332 = n3276 ^ n3272 ;
  assign n3335 = n3331 & n3332 ;
  assign n3340 = n3336 ^ n3335 ;
  assign n3345 = n3343 ^ n3340 ;
  assign n3346 = n3345 ^ n3329 ;
  assign n3298 = n3269 ^ n3265 ;
  assign n3299 = n3270 ^ n3266 ;
  assign n3301 = n3298 & n3299 ;
  assign n3296 = n3267 ^ n3263 ;
  assign n3297 = n3268 ^ n3264 ;
  assign n3300 = n3296 & n3297 ;
  assign n3305 = n3301 ^ n3300 ;
  assign n3310 = n3308 ^ n3305 ;
  assign n3311 = n3310 ^ n3294 ;
  assign n3397 = n3346 ^ n3311 ;
  assign n3419 = n3409 ^ n3397 ;
  assign n3420 = n3419 ^ n3253 ;
  assign n4350 = n3851 ^ n3420 ;
  assign n4440 = n4398 ^ n4350 ;
  assign n4441 = n4440 ^ n2894 ;
  assign n3768 = n3764 ^ n3762 ;
  assign n3769 = n3765 ^ n3763 ;
  assign n3770 = n3768 & n3769 ;
  assign n3772 = n3771 ^ n3770 ;
  assign n3773 = n3772 ^ n3767 ;
  assign n3778 = n3775 ^ n3773 ;
  assign n3761 = n3760 ^ n3758 ;
  assign n3779 = n3778 ^ n3761 ;
  assign n3733 = n3729 ^ n3727 ;
  assign n3734 = n3730 ^ n3728 ;
  assign n3735 = n3733 & n3734 ;
  assign n3737 = n3736 ^ n3735 ;
  assign n3738 = n3737 ^ n3732 ;
  assign n3743 = n3740 ^ n3738 ;
  assign n3726 = n3725 ^ n3723 ;
  assign n3744 = n3743 ^ n3726 ;
  assign n3829 = n3779 ^ n3744 ;
  assign n3852 = n3841 ^ n3829 ;
  assign n3853 = n3852 ^ n3686 ;
  assign n3337 = n3333 ^ n3331 ;
  assign n3338 = n3334 ^ n3332 ;
  assign n3339 = n3337 & n3338 ;
  assign n3341 = n3340 ^ n3339 ;
  assign n3342 = n3341 ^ n3336 ;
  assign n3347 = n3344 ^ n3342 ;
  assign n3330 = n3329 ^ n3327 ;
  assign n3348 = n3347 ^ n3330 ;
  assign n3302 = n3298 ^ n3296 ;
  assign n3303 = n3299 ^ n3297 ;
  assign n3304 = n3302 & n3303 ;
  assign n3306 = n3305 ^ n3304 ;
  assign n3307 = n3306 ^ n3301 ;
  assign n3312 = n3309 ^ n3307 ;
  assign n3295 = n3294 ^ n3292 ;
  assign n3313 = n3312 ^ n3295 ;
  assign n3398 = n3348 ^ n3313 ;
  assign n3421 = n3410 ^ n3398 ;
  assign n3422 = n3421 ^ n3255 ;
  assign n4351 = n3853 ^ n3422 ;
  assign n4442 = n4399 ^ n4351 ;
  assign n4443 = n4442 ^ n2896 ;
  assign n3789 = n3708 ^ n3700 ;
  assign n3790 = n3709 ^ n3701 ;
  assign n3800 = n3789 & n3790 ;
  assign n3787 = n3706 ^ n3698 ;
  assign n3788 = n3707 ^ n3699 ;
  assign n3799 = n3787 & n3788 ;
  assign n3804 = n3800 ^ n3799 ;
  assign n3785 = n3704 ^ n3696 ;
  assign n3786 = n3705 ^ n3697 ;
  assign n3792 = n3785 & n3786 ;
  assign n3783 = n3702 ^ n3694 ;
  assign n3784 = n3703 ^ n3695 ;
  assign n3791 = n3783 & n3784 ;
  assign n3796 = n3792 ^ n3791 ;
  assign n3820 = n3804 ^ n3796 ;
  assign n3830 = n3826 ^ n3820 ;
  assign n3831 = n3830 ^ n3777 ;
  assign n3854 = n3842 ^ n3831 ;
  assign n3690 = n3684 ^ n3675 ;
  assign n3855 = n3854 ^ n3690 ;
  assign n3358 = n3277 ^ n3269 ;
  assign n3359 = n3278 ^ n3270 ;
  assign n3369 = n3358 & n3359 ;
  assign n3356 = n3275 ^ n3267 ;
  assign n3357 = n3276 ^ n3268 ;
  assign n3368 = n3356 & n3357 ;
  assign n3373 = n3369 ^ n3368 ;
  assign n3354 = n3273 ^ n3265 ;
  assign n3355 = n3274 ^ n3266 ;
  assign n3361 = n3354 & n3355 ;
  assign n3352 = n3271 ^ n3263 ;
  assign n3353 = n3272 ^ n3264 ;
  assign n3360 = n3352 & n3353 ;
  assign n3365 = n3361 ^ n3360 ;
  assign n3389 = n3373 ^ n3365 ;
  assign n3399 = n3395 ^ n3389 ;
  assign n3400 = n3399 ^ n3346 ;
  assign n3423 = n3411 ^ n3400 ;
  assign n3259 = n3253 ^ n3244 ;
  assign n3424 = n3423 ^ n3259 ;
  assign n4352 = n3855 ^ n3424 ;
  assign n4444 = n4400 ^ n4352 ;
  assign n4445 = n4444 ^ n2898 ;
  assign n3801 = n3789 ^ n3787 ;
  assign n3802 = n3790 ^ n3788 ;
  assign n3803 = n3801 & n3802 ;
  assign n3805 = n3804 ^ n3803 ;
  assign n3806 = n3805 ^ n3800 ;
  assign n3793 = n3785 ^ n3783 ;
  assign n3794 = n3786 ^ n3784 ;
  assign n3795 = n3793 & n3794 ;
  assign n3797 = n3796 ^ n3795 ;
  assign n3798 = n3797 ^ n3792 ;
  assign n3821 = n3806 ^ n3798 ;
  assign n3832 = n3827 ^ n3821 ;
  assign n3833 = n3832 ^ n3779 ;
  assign n3856 = n3843 ^ n3833 ;
  assign n3691 = n3686 ^ n3676 ;
  assign n3857 = n3856 ^ n3691 ;
  assign n3370 = n3358 ^ n3356 ;
  assign n3371 = n3359 ^ n3357 ;
  assign n3372 = n3370 & n3371 ;
  assign n3374 = n3373 ^ n3372 ;
  assign n3375 = n3374 ^ n3369 ;
  assign n3362 = n3354 ^ n3352 ;
  assign n3363 = n3355 ^ n3353 ;
  assign n3364 = n3362 & n3363 ;
  assign n3366 = n3365 ^ n3364 ;
  assign n3367 = n3366 ^ n3361 ;
  assign n3390 = n3375 ^ n3367 ;
  assign n3401 = n3396 ^ n3390 ;
  assign n3402 = n3401 ^ n3348 ;
  assign n3425 = n3412 ^ n3402 ;
  assign n3260 = n3255 ^ n3245 ;
  assign n3426 = n3425 ^ n3260 ;
  assign n4353 = n3857 ^ n3426 ;
  assign n4446 = n4401 ^ n4353 ;
  assign n4447 = n4446 ^ n2900 ;
  assign n3810 = n3789 ^ n3785 ;
  assign n3811 = n3790 ^ n3786 ;
  assign n3813 = n3810 & n3811 ;
  assign n3808 = n3787 ^ n3783 ;
  assign n3809 = n3788 ^ n3784 ;
  assign n3812 = n3808 & n3809 ;
  assign n3817 = n3813 ^ n3812 ;
  assign n3822 = n3820 ^ n3817 ;
  assign n3823 = n3822 ^ n3806 ;
  assign n3834 = n3828 ^ n3823 ;
  assign n3781 = n3779 ^ n3774 ;
  assign n3835 = n3834 ^ n3781 ;
  assign n3858 = n3844 ^ n3835 ;
  assign n3688 = n3686 ^ n3680 ;
  assign n3692 = n3688 ^ n3677 ;
  assign n3859 = n3858 ^ n3692 ;
  assign n3379 = n3358 ^ n3354 ;
  assign n3380 = n3359 ^ n3355 ;
  assign n3382 = n3379 & n3380 ;
  assign n3377 = n3356 ^ n3352 ;
  assign n3378 = n3357 ^ n3353 ;
  assign n3381 = n3377 & n3378 ;
  assign n3386 = n3382 ^ n3381 ;
  assign n3391 = n3389 ^ n3386 ;
  assign n3392 = n3391 ^ n3375 ;
  assign n3403 = n3397 ^ n3392 ;
  assign n3350 = n3348 ^ n3343 ;
  assign n3404 = n3403 ^ n3350 ;
  assign n3427 = n3413 ^ n3404 ;
  assign n3257 = n3255 ^ n3249 ;
  assign n3261 = n3257 ^ n3246 ;
  assign n3428 = n3427 ^ n3261 ;
  assign n4354 = n3859 ^ n3428 ;
  assign n4448 = n4402 ^ n4354 ;
  assign n4449 = n4448 ^ n2902 ;
  assign n3814 = n3810 ^ n3808 ;
  assign n3815 = n3811 ^ n3809 ;
  assign n3816 = n3814 & n3815 ;
  assign n3818 = n3817 ^ n3816 ;
  assign n3819 = n3818 ^ n3813 ;
  assign n3824 = n3821 ^ n3819 ;
  assign n3807 = n3806 ^ n3804 ;
  assign n3825 = n3824 ^ n3807 ;
  assign n3836 = n3829 ^ n3825 ;
  assign n3780 = n3779 ^ n3777 ;
  assign n3782 = n3780 ^ n3775 ;
  assign n3837 = n3836 ^ n3782 ;
  assign n3860 = n3845 ^ n3837 ;
  assign n3687 = n3686 ^ n3684 ;
  assign n3689 = n3687 ^ n3682 ;
  assign n3693 = n3689 ^ n3678 ;
  assign n3861 = n3860 ^ n3693 ;
  assign n3383 = n3379 ^ n3377 ;
  assign n3384 = n3380 ^ n3378 ;
  assign n3385 = n3383 & n3384 ;
  assign n3387 = n3386 ^ n3385 ;
  assign n3388 = n3387 ^ n3382 ;
  assign n3393 = n3390 ^ n3388 ;
  assign n3376 = n3375 ^ n3373 ;
  assign n3394 = n3393 ^ n3376 ;
  assign n3405 = n3398 ^ n3394 ;
  assign n3349 = n3348 ^ n3346 ;
  assign n3351 = n3349 ^ n3344 ;
  assign n3406 = n3405 ^ n3351 ;
  assign n3429 = n3414 ^ n3406 ;
  assign n3256 = n3255 ^ n3253 ;
  assign n3258 = n3256 ^ n3251 ;
  assign n3262 = n3258 ^ n3247 ;
  assign n3430 = n3429 ^ n3262 ;
  assign n4355 = n3861 ^ n3430 ;
  assign n4450 = n4403 ^ n4355 ;
  assign n4451 = n4450 ^ n2904 ;
  assign n3907 = n2998 ^ n2966 ;
  assign n3908 = n2999 ^ n2967 ;
  assign n4081 = n3907 & n3908 ;
  assign n3905 = n2996 ^ n2964 ;
  assign n3906 = n2997 ^ n2965 ;
  assign n4080 = n3905 & n3906 ;
  assign n4085 = n4081 ^ n4080 ;
  assign n3903 = n2994 ^ n2962 ;
  assign n3904 = n2995 ^ n2963 ;
  assign n4073 = n3903 & n3904 ;
  assign n3901 = n2992 ^ n2960 ;
  assign n3902 = n2993 ^ n2961 ;
  assign n4072 = n3901 & n3902 ;
  assign n4077 = n4073 ^ n4072 ;
  assign n4101 = n4085 ^ n4077 ;
  assign n3899 = n2990 ^ n2958 ;
  assign n3900 = n2991 ^ n2959 ;
  assign n4046 = n3899 & n3900 ;
  assign n3897 = n2988 ^ n2956 ;
  assign n3898 = n2989 ^ n2957 ;
  assign n4045 = n3897 & n3898 ;
  assign n4050 = n4046 ^ n4045 ;
  assign n3895 = n2986 ^ n2954 ;
  assign n3896 = n2987 ^ n2955 ;
  assign n4038 = n3895 & n3896 ;
  assign n3893 = n2984 ^ n2952 ;
  assign n3894 = n2985 ^ n2953 ;
  assign n4037 = n3893 & n3894 ;
  assign n4042 = n4038 ^ n4037 ;
  assign n4066 = n4050 ^ n4042 ;
  assign n4153 = n4101 ^ n4066 ;
  assign n3891 = n2982 ^ n2950 ;
  assign n3892 = n2983 ^ n2951 ;
  assign n3953 = n3891 & n3892 ;
  assign n3889 = n2980 ^ n2948 ;
  assign n3890 = n2981 ^ n2949 ;
  assign n3952 = n3889 & n3890 ;
  assign n3957 = n3953 ^ n3952 ;
  assign n3887 = n2978 ^ n2946 ;
  assign n3888 = n2979 ^ n2947 ;
  assign n3945 = n3887 & n3888 ;
  assign n3885 = n2976 ^ n2944 ;
  assign n3886 = n2977 ^ n2945 ;
  assign n3944 = n3885 & n3886 ;
  assign n3949 = n3945 ^ n3944 ;
  assign n3973 = n3957 ^ n3949 ;
  assign n3883 = n2974 ^ n2942 ;
  assign n3884 = n2975 ^ n2943 ;
  assign n3918 = n3883 & n3884 ;
  assign n3881 = n2972 ^ n2940 ;
  assign n3882 = n2973 ^ n2941 ;
  assign n3917 = n3881 & n3882 ;
  assign n3922 = n3918 ^ n3917 ;
  assign n3879 = n2970 ^ n2938 ;
  assign n3880 = n2971 ^ n2939 ;
  assign n3910 = n3879 & n3880 ;
  assign n3877 = n2968 ^ n2936 ;
  assign n3878 = n2969 ^ n2937 ;
  assign n3909 = n3877 & n3878 ;
  assign n3914 = n3910 ^ n3909 ;
  assign n3938 = n3922 ^ n3914 ;
  assign n4025 = n3973 ^ n3938 ;
  assign n4316 = n4153 ^ n4025 ;
  assign n4356 = n4340 ^ n4316 ;
  assign n4357 = n4356 ^ n3847 ;
  assign n4452 = n4404 ^ n4357 ;
  assign n2920 = n2890 ^ n2857 ;
  assign n4453 = n4452 ^ n2920 ;
  assign n4082 = n3907 ^ n3905 ;
  assign n4083 = n3908 ^ n3906 ;
  assign n4084 = n4082 & n4083 ;
  assign n4086 = n4085 ^ n4084 ;
  assign n4087 = n4086 ^ n4081 ;
  assign n4074 = n3903 ^ n3901 ;
  assign n4075 = n3904 ^ n3902 ;
  assign n4076 = n4074 & n4075 ;
  assign n4078 = n4077 ^ n4076 ;
  assign n4079 = n4078 ^ n4073 ;
  assign n4102 = n4087 ^ n4079 ;
  assign n4047 = n3899 ^ n3897 ;
  assign n4048 = n3900 ^ n3898 ;
  assign n4049 = n4047 & n4048 ;
  assign n4051 = n4050 ^ n4049 ;
  assign n4052 = n4051 ^ n4046 ;
  assign n4039 = n3895 ^ n3893 ;
  assign n4040 = n3896 ^ n3894 ;
  assign n4041 = n4039 & n4040 ;
  assign n4043 = n4042 ^ n4041 ;
  assign n4044 = n4043 ^ n4038 ;
  assign n4067 = n4052 ^ n4044 ;
  assign n4154 = n4102 ^ n4067 ;
  assign n3954 = n3891 ^ n3889 ;
  assign n3955 = n3892 ^ n3890 ;
  assign n3956 = n3954 & n3955 ;
  assign n3958 = n3957 ^ n3956 ;
  assign n3959 = n3958 ^ n3953 ;
  assign n3946 = n3887 ^ n3885 ;
  assign n3947 = n3888 ^ n3886 ;
  assign n3948 = n3946 & n3947 ;
  assign n3950 = n3949 ^ n3948 ;
  assign n3951 = n3950 ^ n3945 ;
  assign n3974 = n3959 ^ n3951 ;
  assign n3919 = n3883 ^ n3881 ;
  assign n3920 = n3884 ^ n3882 ;
  assign n3921 = n3919 & n3920 ;
  assign n3923 = n3922 ^ n3921 ;
  assign n3924 = n3923 ^ n3918 ;
  assign n3911 = n3879 ^ n3877 ;
  assign n3912 = n3880 ^ n3878 ;
  assign n3913 = n3911 & n3912 ;
  assign n3915 = n3914 ^ n3913 ;
  assign n3916 = n3915 ^ n3910 ;
  assign n3939 = n3924 ^ n3916 ;
  assign n4026 = n3974 ^ n3939 ;
  assign n4317 = n4154 ^ n4026 ;
  assign n4358 = n4341 ^ n4317 ;
  assign n4359 = n4358 ^ n3849 ;
  assign n4454 = n4405 ^ n4359 ;
  assign n2921 = n2892 ^ n2858 ;
  assign n4455 = n4454 ^ n2921 ;
  assign n4091 = n3907 ^ n3903 ;
  assign n4092 = n3908 ^ n3904 ;
  assign n4094 = n4091 & n4092 ;
  assign n4089 = n3905 ^ n3901 ;
  assign n4090 = n3906 ^ n3902 ;
  assign n4093 = n4089 & n4090 ;
  assign n4098 = n4094 ^ n4093 ;
  assign n4103 = n4101 ^ n4098 ;
  assign n4104 = n4103 ^ n4087 ;
  assign n4056 = n3899 ^ n3895 ;
  assign n4057 = n3900 ^ n3896 ;
  assign n4059 = n4056 & n4057 ;
  assign n4054 = n3897 ^ n3893 ;
  assign n4055 = n3898 ^ n3894 ;
  assign n4058 = n4054 & n4055 ;
  assign n4063 = n4059 ^ n4058 ;
  assign n4068 = n4066 ^ n4063 ;
  assign n4069 = n4068 ^ n4052 ;
  assign n4155 = n4104 ^ n4069 ;
  assign n3963 = n3891 ^ n3887 ;
  assign n3964 = n3892 ^ n3888 ;
  assign n3966 = n3963 & n3964 ;
  assign n3961 = n3889 ^ n3885 ;
  assign n3962 = n3890 ^ n3886 ;
  assign n3965 = n3961 & n3962 ;
  assign n3970 = n3966 ^ n3965 ;
  assign n3975 = n3973 ^ n3970 ;
  assign n3976 = n3975 ^ n3959 ;
  assign n3928 = n3883 ^ n3879 ;
  assign n3929 = n3884 ^ n3880 ;
  assign n3931 = n3928 & n3929 ;
  assign n3926 = n3881 ^ n3877 ;
  assign n3927 = n3882 ^ n3878 ;
  assign n3930 = n3926 & n3927 ;
  assign n3935 = n3931 ^ n3930 ;
  assign n3940 = n3938 ^ n3935 ;
  assign n3941 = n3940 ^ n3924 ;
  assign n4027 = n3976 ^ n3941 ;
  assign n4318 = n4155 ^ n4027 ;
  assign n4360 = n4342 ^ n4318 ;
  assign n4361 = n4360 ^ n3851 ;
  assign n4456 = n4406 ^ n4361 ;
  assign n2922 = n2894 ^ n2859 ;
  assign n4457 = n4456 ^ n2922 ;
  assign n4095 = n4091 ^ n4089 ;
  assign n4096 = n4092 ^ n4090 ;
  assign n4097 = n4095 & n4096 ;
  assign n4099 = n4098 ^ n4097 ;
  assign n4100 = n4099 ^ n4094 ;
  assign n4105 = n4102 ^ n4100 ;
  assign n4088 = n4087 ^ n4085 ;
  assign n4106 = n4105 ^ n4088 ;
  assign n4060 = n4056 ^ n4054 ;
  assign n4061 = n4057 ^ n4055 ;
  assign n4062 = n4060 & n4061 ;
  assign n4064 = n4063 ^ n4062 ;
  assign n4065 = n4064 ^ n4059 ;
  assign n4070 = n4067 ^ n4065 ;
  assign n4053 = n4052 ^ n4050 ;
  assign n4071 = n4070 ^ n4053 ;
  assign n4156 = n4106 ^ n4071 ;
  assign n3967 = n3963 ^ n3961 ;
  assign n3968 = n3964 ^ n3962 ;
  assign n3969 = n3967 & n3968 ;
  assign n3971 = n3970 ^ n3969 ;
  assign n3972 = n3971 ^ n3966 ;
  assign n3977 = n3974 ^ n3972 ;
  assign n3960 = n3959 ^ n3957 ;
  assign n3978 = n3977 ^ n3960 ;
  assign n3932 = n3928 ^ n3926 ;
  assign n3933 = n3929 ^ n3927 ;
  assign n3934 = n3932 & n3933 ;
  assign n3936 = n3935 ^ n3934 ;
  assign n3937 = n3936 ^ n3931 ;
  assign n3942 = n3939 ^ n3937 ;
  assign n3925 = n3924 ^ n3922 ;
  assign n3943 = n3942 ^ n3925 ;
  assign n4028 = n3978 ^ n3943 ;
  assign n4319 = n4156 ^ n4028 ;
  assign n4362 = n4343 ^ n4319 ;
  assign n4363 = n4362 ^ n3853 ;
  assign n4458 = n4407 ^ n4363 ;
  assign n2923 = n2896 ^ n2860 ;
  assign n4459 = n4458 ^ n2923 ;
  assign n4116 = n3907 ^ n3899 ;
  assign n4117 = n3908 ^ n3900 ;
  assign n4127 = n4116 & n4117 ;
  assign n4114 = n3905 ^ n3897 ;
  assign n4115 = n3906 ^ n3898 ;
  assign n4126 = n4114 & n4115 ;
  assign n4131 = n4127 ^ n4126 ;
  assign n4112 = n3903 ^ n3895 ;
  assign n4113 = n3904 ^ n3896 ;
  assign n4119 = n4112 & n4113 ;
  assign n4110 = n3901 ^ n3893 ;
  assign n4111 = n3902 ^ n3894 ;
  assign n4118 = n4110 & n4111 ;
  assign n4123 = n4119 ^ n4118 ;
  assign n4147 = n4131 ^ n4123 ;
  assign n4157 = n4153 ^ n4147 ;
  assign n4158 = n4157 ^ n4104 ;
  assign n3988 = n3891 ^ n3883 ;
  assign n3989 = n3892 ^ n3884 ;
  assign n3999 = n3988 & n3989 ;
  assign n3986 = n3889 ^ n3881 ;
  assign n3987 = n3890 ^ n3882 ;
  assign n3998 = n3986 & n3987 ;
  assign n4003 = n3999 ^ n3998 ;
  assign n3984 = n3887 ^ n3879 ;
  assign n3985 = n3888 ^ n3880 ;
  assign n3991 = n3984 & n3985 ;
  assign n3982 = n3885 ^ n3877 ;
  assign n3983 = n3886 ^ n3878 ;
  assign n3990 = n3982 & n3983 ;
  assign n3995 = n3991 ^ n3990 ;
  assign n4019 = n4003 ^ n3995 ;
  assign n4029 = n4025 ^ n4019 ;
  assign n4030 = n4029 ^ n3976 ;
  assign n4320 = n4158 ^ n4030 ;
  assign n4364 = n4344 ^ n4320 ;
  assign n4365 = n4364 ^ n3855 ;
  assign n4460 = n4408 ^ n4365 ;
  assign n2924 = n2898 ^ n2861 ;
  assign n4461 = n4460 ^ n2924 ;
  assign n4128 = n4116 ^ n4114 ;
  assign n4129 = n4117 ^ n4115 ;
  assign n4130 = n4128 & n4129 ;
  assign n4132 = n4131 ^ n4130 ;
  assign n4133 = n4132 ^ n4127 ;
  assign n4120 = n4112 ^ n4110 ;
  assign n4121 = n4113 ^ n4111 ;
  assign n4122 = n4120 & n4121 ;
  assign n4124 = n4123 ^ n4122 ;
  assign n4125 = n4124 ^ n4119 ;
  assign n4148 = n4133 ^ n4125 ;
  assign n4159 = n4154 ^ n4148 ;
  assign n4160 = n4159 ^ n4106 ;
  assign n4000 = n3988 ^ n3986 ;
  assign n4001 = n3989 ^ n3987 ;
  assign n4002 = n4000 & n4001 ;
  assign n4004 = n4003 ^ n4002 ;
  assign n4005 = n4004 ^ n3999 ;
  assign n3992 = n3984 ^ n3982 ;
  assign n3993 = n3985 ^ n3983 ;
  assign n3994 = n3992 & n3993 ;
  assign n3996 = n3995 ^ n3994 ;
  assign n3997 = n3996 ^ n3991 ;
  assign n4020 = n4005 ^ n3997 ;
  assign n4031 = n4026 ^ n4020 ;
  assign n4032 = n4031 ^ n3978 ;
  assign n4321 = n4160 ^ n4032 ;
  assign n4366 = n4345 ^ n4321 ;
  assign n4367 = n4366 ^ n3857 ;
  assign n4462 = n4409 ^ n4367 ;
  assign n2925 = n2900 ^ n2862 ;
  assign n4463 = n4462 ^ n2925 ;
  assign n4137 = n4116 ^ n4112 ;
  assign n4138 = n4117 ^ n4113 ;
  assign n4140 = n4137 & n4138 ;
  assign n4135 = n4114 ^ n4110 ;
  assign n4136 = n4115 ^ n4111 ;
  assign n4139 = n4135 & n4136 ;
  assign n4144 = n4140 ^ n4139 ;
  assign n4149 = n4147 ^ n4144 ;
  assign n4150 = n4149 ^ n4133 ;
  assign n4161 = n4155 ^ n4150 ;
  assign n4108 = n4106 ^ n4101 ;
  assign n4162 = n4161 ^ n4108 ;
  assign n4009 = n3988 ^ n3984 ;
  assign n4010 = n3989 ^ n3985 ;
  assign n4012 = n4009 & n4010 ;
  assign n4007 = n3986 ^ n3982 ;
  assign n4008 = n3987 ^ n3983 ;
  assign n4011 = n4007 & n4008 ;
  assign n4016 = n4012 ^ n4011 ;
  assign n4021 = n4019 ^ n4016 ;
  assign n4022 = n4021 ^ n4005 ;
  assign n4033 = n4027 ^ n4022 ;
  assign n3980 = n3978 ^ n3973 ;
  assign n4034 = n4033 ^ n3980 ;
  assign n4322 = n4162 ^ n4034 ;
  assign n4368 = n4346 ^ n4322 ;
  assign n4369 = n4368 ^ n3859 ;
  assign n4464 = n4410 ^ n4369 ;
  assign n2926 = n2902 ^ n2863 ;
  assign n4465 = n4464 ^ n2926 ;
  assign n4141 = n4137 ^ n4135 ;
  assign n4142 = n4138 ^ n4136 ;
  assign n4143 = n4141 & n4142 ;
  assign n4145 = n4144 ^ n4143 ;
  assign n4146 = n4145 ^ n4140 ;
  assign n4151 = n4148 ^ n4146 ;
  assign n4134 = n4133 ^ n4131 ;
  assign n4152 = n4151 ^ n4134 ;
  assign n4163 = n4156 ^ n4152 ;
  assign n4107 = n4106 ^ n4104 ;
  assign n4109 = n4107 ^ n4102 ;
  assign n4164 = n4163 ^ n4109 ;
  assign n4013 = n4009 ^ n4007 ;
  assign n4014 = n4010 ^ n4008 ;
  assign n4015 = n4013 & n4014 ;
  assign n4017 = n4016 ^ n4015 ;
  assign n4018 = n4017 ^ n4012 ;
  assign n4023 = n4020 ^ n4018 ;
  assign n4006 = n4005 ^ n4003 ;
  assign n4024 = n4023 ^ n4006 ;
  assign n4035 = n4028 ^ n4024 ;
  assign n3979 = n3978 ^ n3976 ;
  assign n3981 = n3979 ^ n3974 ;
  assign n4036 = n4035 ^ n3981 ;
  assign n4323 = n4164 ^ n4036 ;
  assign n4370 = n4347 ^ n4323 ;
  assign n4371 = n4370 ^ n3861 ;
  assign n4466 = n4411 ^ n4371 ;
  assign n2927 = n2904 ^ n2864 ;
  assign n4467 = n4466 ^ n2927 ;
  assign n4186 = n3907 ^ n3891 ;
  assign n4187 = n3908 ^ n3892 ;
  assign n4232 = n4186 & n4187 ;
  assign n4184 = n3905 ^ n3889 ;
  assign n4185 = n3906 ^ n3890 ;
  assign n4231 = n4184 & n4185 ;
  assign n4236 = n4232 ^ n4231 ;
  assign n4182 = n3903 ^ n3887 ;
  assign n4183 = n3904 ^ n3888 ;
  assign n4224 = n4182 & n4183 ;
  assign n4180 = n3901 ^ n3885 ;
  assign n4181 = n3902 ^ n3886 ;
  assign n4223 = n4180 & n4181 ;
  assign n4228 = n4224 ^ n4223 ;
  assign n4252 = n4236 ^ n4228 ;
  assign n4178 = n3899 ^ n3883 ;
  assign n4179 = n3900 ^ n3884 ;
  assign n4197 = n4178 & n4179 ;
  assign n4176 = n3897 ^ n3881 ;
  assign n4177 = n3898 ^ n3882 ;
  assign n4196 = n4176 & n4177 ;
  assign n4201 = n4197 ^ n4196 ;
  assign n4174 = n3895 ^ n3879 ;
  assign n4175 = n3896 ^ n3880 ;
  assign n4189 = n4174 & n4175 ;
  assign n4172 = n3893 ^ n3877 ;
  assign n4173 = n3894 ^ n3878 ;
  assign n4188 = n4172 & n4173 ;
  assign n4193 = n4189 ^ n4188 ;
  assign n4217 = n4201 ^ n4193 ;
  assign n4304 = n4252 ^ n4217 ;
  assign n4324 = n4316 ^ n4304 ;
  assign n4325 = n4324 ^ n4158 ;
  assign n4372 = n4348 ^ n4325 ;
  assign n3869 = n3855 ^ n3838 ;
  assign n4373 = n4372 ^ n3869 ;
  assign n4468 = n4412 ^ n4373 ;
  assign n2912 = n2898 ^ n2874 ;
  assign n2928 = n2912 ^ n2865 ;
  assign n4469 = n4468 ^ n2928 ;
  assign n4233 = n4186 ^ n4184 ;
  assign n4234 = n4187 ^ n4185 ;
  assign n4235 = n4233 & n4234 ;
  assign n4237 = n4236 ^ n4235 ;
  assign n4238 = n4237 ^ n4232 ;
  assign n4225 = n4182 ^ n4180 ;
  assign n4226 = n4183 ^ n4181 ;
  assign n4227 = n4225 & n4226 ;
  assign n4229 = n4228 ^ n4227 ;
  assign n4230 = n4229 ^ n4224 ;
  assign n4253 = n4238 ^ n4230 ;
  assign n4198 = n4178 ^ n4176 ;
  assign n4199 = n4179 ^ n4177 ;
  assign n4200 = n4198 & n4199 ;
  assign n4202 = n4201 ^ n4200 ;
  assign n4203 = n4202 ^ n4197 ;
  assign n4190 = n4174 ^ n4172 ;
  assign n4191 = n4175 ^ n4173 ;
  assign n4192 = n4190 & n4191 ;
  assign n4194 = n4193 ^ n4192 ;
  assign n4195 = n4194 ^ n4189 ;
  assign n4218 = n4203 ^ n4195 ;
  assign n4305 = n4253 ^ n4218 ;
  assign n4326 = n4317 ^ n4305 ;
  assign n4327 = n4326 ^ n4160 ;
  assign n4374 = n4349 ^ n4327 ;
  assign n3870 = n3857 ^ n3839 ;
  assign n4375 = n4374 ^ n3870 ;
  assign n4470 = n4413 ^ n4375 ;
  assign n2913 = n2900 ^ n2876 ;
  assign n2929 = n2913 ^ n2866 ;
  assign n4471 = n4470 ^ n2929 ;
  assign n4242 = n4186 ^ n4182 ;
  assign n4243 = n4187 ^ n4183 ;
  assign n4245 = n4242 & n4243 ;
  assign n4240 = n4184 ^ n4180 ;
  assign n4241 = n4185 ^ n4181 ;
  assign n4244 = n4240 & n4241 ;
  assign n4249 = n4245 ^ n4244 ;
  assign n4254 = n4252 ^ n4249 ;
  assign n4255 = n4254 ^ n4238 ;
  assign n4207 = n4178 ^ n4174 ;
  assign n4208 = n4179 ^ n4175 ;
  assign n4210 = n4207 & n4208 ;
  assign n4205 = n4176 ^ n4172 ;
  assign n4206 = n4177 ^ n4173 ;
  assign n4209 = n4205 & n4206 ;
  assign n4214 = n4210 ^ n4209 ;
  assign n4219 = n4217 ^ n4214 ;
  assign n4220 = n4219 ^ n4203 ;
  assign n4306 = n4255 ^ n4220 ;
  assign n4328 = n4318 ^ n4306 ;
  assign n4329 = n4328 ^ n4162 ;
  assign n4376 = n4350 ^ n4329 ;
  assign n3871 = n3859 ^ n3840 ;
  assign n4377 = n4376 ^ n3871 ;
  assign n4472 = n4414 ^ n4377 ;
  assign n2914 = n2902 ^ n2878 ;
  assign n2930 = n2914 ^ n2867 ;
  assign n4473 = n4472 ^ n2930 ;
  assign n4246 = n4242 ^ n4240 ;
  assign n4247 = n4243 ^ n4241 ;
  assign n4248 = n4246 & n4247 ;
  assign n4250 = n4249 ^ n4248 ;
  assign n4251 = n4250 ^ n4245 ;
  assign n4256 = n4253 ^ n4251 ;
  assign n4239 = n4238 ^ n4236 ;
  assign n4257 = n4256 ^ n4239 ;
  assign n4211 = n4207 ^ n4205 ;
  assign n4212 = n4208 ^ n4206 ;
  assign n4213 = n4211 & n4212 ;
  assign n4215 = n4214 ^ n4213 ;
  assign n4216 = n4215 ^ n4210 ;
  assign n4221 = n4218 ^ n4216 ;
  assign n4204 = n4203 ^ n4201 ;
  assign n4222 = n4221 ^ n4204 ;
  assign n4307 = n4257 ^ n4222 ;
  assign n4330 = n4319 ^ n4307 ;
  assign n4331 = n4330 ^ n4164 ;
  assign n4378 = n4351 ^ n4331 ;
  assign n3872 = n3861 ^ n3841 ;
  assign n4379 = n4378 ^ n3872 ;
  assign n4474 = n4415 ^ n4379 ;
  assign n2915 = n2904 ^ n2880 ;
  assign n2931 = n2915 ^ n2868 ;
  assign n4475 = n4474 ^ n2931 ;
  assign n4267 = n4186 ^ n4178 ;
  assign n4268 = n4187 ^ n4179 ;
  assign n4278 = n4267 & n4268 ;
  assign n4265 = n4184 ^ n4176 ;
  assign n4266 = n4185 ^ n4177 ;
  assign n4277 = n4265 & n4266 ;
  assign n4282 = n4278 ^ n4277 ;
  assign n4263 = n4182 ^ n4174 ;
  assign n4264 = n4183 ^ n4175 ;
  assign n4270 = n4263 & n4264 ;
  assign n4261 = n4180 ^ n4172 ;
  assign n4262 = n4181 ^ n4173 ;
  assign n4269 = n4261 & n4262 ;
  assign n4274 = n4270 ^ n4269 ;
  assign n4298 = n4282 ^ n4274 ;
  assign n4308 = n4304 ^ n4298 ;
  assign n4309 = n4308 ^ n4255 ;
  assign n4332 = n4320 ^ n4309 ;
  assign n4168 = n4162 ^ n4153 ;
  assign n4333 = n4332 ^ n4168 ;
  assign n4380 = n4352 ^ n4333 ;
  assign n3865 = n3859 ^ n3847 ;
  assign n3873 = n3865 ^ n3842 ;
  assign n4381 = n4380 ^ n3873 ;
  assign n4476 = n4416 ^ n4381 ;
  assign n2908 = n2902 ^ n2890 ;
  assign n2916 = n2908 ^ n2882 ;
  assign n2932 = n2916 ^ n2869 ;
  assign n4477 = n4476 ^ n2932 ;
  assign n4279 = n4267 ^ n4265 ;
  assign n4280 = n4268 ^ n4266 ;
  assign n4281 = n4279 & n4280 ;
  assign n4283 = n4282 ^ n4281 ;
  assign n4284 = n4283 ^ n4278 ;
  assign n4271 = n4263 ^ n4261 ;
  assign n4272 = n4264 ^ n4262 ;
  assign n4273 = n4271 & n4272 ;
  assign n4275 = n4274 ^ n4273 ;
  assign n4276 = n4275 ^ n4270 ;
  assign n4299 = n4284 ^ n4276 ;
  assign n4310 = n4305 ^ n4299 ;
  assign n4311 = n4310 ^ n4257 ;
  assign n4334 = n4321 ^ n4311 ;
  assign n4169 = n4164 ^ n4154 ;
  assign n4335 = n4334 ^ n4169 ;
  assign n4382 = n4353 ^ n4335 ;
  assign n3866 = n3861 ^ n3849 ;
  assign n3874 = n3866 ^ n3843 ;
  assign n4383 = n4382 ^ n3874 ;
  assign n4478 = n4417 ^ n4383 ;
  assign n2909 = n2904 ^ n2892 ;
  assign n2917 = n2909 ^ n2884 ;
  assign n2933 = n2917 ^ n2870 ;
  assign n4479 = n4478 ^ n2933 ;
  assign n4288 = n4267 ^ n4263 ;
  assign n4289 = n4268 ^ n4264 ;
  assign n4291 = n4288 & n4289 ;
  assign n4286 = n4265 ^ n4261 ;
  assign n4287 = n4266 ^ n4262 ;
  assign n4290 = n4286 & n4287 ;
  assign n4295 = n4291 ^ n4290 ;
  assign n4300 = n4298 ^ n4295 ;
  assign n4301 = n4300 ^ n4284 ;
  assign n4312 = n4306 ^ n4301 ;
  assign n4259 = n4257 ^ n4252 ;
  assign n4313 = n4312 ^ n4259 ;
  assign n4336 = n4322 ^ n4313 ;
  assign n4166 = n4164 ^ n4158 ;
  assign n4170 = n4166 ^ n4155 ;
  assign n4337 = n4336 ^ n4170 ;
  assign n4384 = n4354 ^ n4337 ;
  assign n3863 = n3861 ^ n3855 ;
  assign n3867 = n3863 ^ n3851 ;
  assign n3875 = n3867 ^ n3844 ;
  assign n4385 = n4384 ^ n3875 ;
  assign n4480 = n4418 ^ n4385 ;
  assign n2906 = n2904 ^ n2898 ;
  assign n2910 = n2906 ^ n2894 ;
  assign n2918 = n2910 ^ n2886 ;
  assign n2934 = n2918 ^ n2871 ;
  assign n4481 = n4480 ^ n2934 ;
  assign n4292 = n4288 ^ n4286 ;
  assign n4293 = n4289 ^ n4287 ;
  assign n4294 = n4292 & n4293 ;
  assign n4296 = n4295 ^ n4294 ;
  assign n4297 = n4296 ^ n4291 ;
  assign n4302 = n4299 ^ n4297 ;
  assign n4285 = n4284 ^ n4282 ;
  assign n4303 = n4302 ^ n4285 ;
  assign n4314 = n4307 ^ n4303 ;
  assign n4258 = n4257 ^ n4255 ;
  assign n4260 = n4258 ^ n4253 ;
  assign n4315 = n4314 ^ n4260 ;
  assign n4338 = n4323 ^ n4315 ;
  assign n4165 = n4164 ^ n4162 ;
  assign n4167 = n4165 ^ n4160 ;
  assign n4171 = n4167 ^ n4156 ;
  assign n4339 = n4338 ^ n4171 ;
  assign n4386 = n4355 ^ n4339 ;
  assign n3862 = n3861 ^ n3859 ;
  assign n3864 = n3862 ^ n3857 ;
  assign n3868 = n3864 ^ n3853 ;
  assign n3876 = n3868 ^ n3845 ;
  assign n4387 = n4386 ^ n3876 ;
  assign n4482 = n4419 ^ n4387 ;
  assign n2905 = n2904 ^ n2902 ;
  assign n2907 = n2905 ^ n2900 ;
  assign n2911 = n2907 ^ n2896 ;
  assign n2919 = n2911 ^ n2888 ;
  assign n2935 = n2919 ^ n2872 ;
  assign n4483 = n4482 ^ n2935 ;
  assign y0 = n4388 ;
  assign y1 = n4389 ;
  assign y2 = n4390 ;
  assign y3 = n4391 ;
  assign y4 = n4392 ;
  assign y5 = n4393 ;
  assign y6 = n4394 ;
  assign y7 = n4395 ;
  assign y8 = n4396 ;
  assign y9 = n4397 ;
  assign y10 = n4398 ;
  assign y11 = n4399 ;
  assign y12 = n4400 ;
  assign y13 = n4401 ;
  assign y14 = n4402 ;
  assign y15 = n4403 ;
  assign y16 = n4404 ;
  assign y17 = n4405 ;
  assign y18 = n4406 ;
  assign y19 = n4407 ;
  assign y20 = n4408 ;
  assign y21 = n4409 ;
  assign y22 = n4410 ;
  assign y23 = n4411 ;
  assign y24 = n4412 ;
  assign y25 = n4413 ;
  assign y26 = n4414 ;
  assign y27 = n4415 ;
  assign y28 = n4416 ;
  assign y29 = n4417 ;
  assign y30 = n4418 ;
  assign y31 = n4419 ;
  assign y32 = n4421 ;
  assign y33 = n4423 ;
  assign y34 = n4425 ;
  assign y35 = n4427 ;
  assign y36 = n4429 ;
  assign y37 = n4431 ;
  assign y38 = n4433 ;
  assign y39 = n4435 ;
  assign y40 = n4437 ;
  assign y41 = n4439 ;
  assign y42 = n4441 ;
  assign y43 = n4443 ;
  assign y44 = n4445 ;
  assign y45 = n4447 ;
  assign y46 = n4449 ;
  assign y47 = n4451 ;
  assign y48 = n4453 ;
  assign y49 = n4455 ;
  assign y50 = n4457 ;
  assign y51 = n4459 ;
  assign y52 = n4461 ;
  assign y53 = n4463 ;
  assign y54 = n4465 ;
  assign y55 = n4467 ;
  assign y56 = n4469 ;
  assign y57 = n4471 ;
  assign y58 = n4473 ;
  assign y59 = n4475 ;
  assign y60 = n4477 ;
  assign y61 = n4479 ;
  assign y62 = n4481 ;
  assign y63 = n4483 ;
endmodule
